module rs_latch_new(
       input top_in_n, 
       input top_in_p, 
       input VDD, 
       input VSS, 
       output top_out_n, 
       output top_out_p 
);

endmodule


