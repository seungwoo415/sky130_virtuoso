VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO DigitalLDOLogic
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DigitalLDOLogic 0 0 ;
  SIZE 200 BY 60 ;
  SYMMETRY X Y ;
  SITE unithd ;
  PIN clk
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 170.185 22.245 170.515 22.615 ;
        RECT 133.385 22.245 133.715 22.615 ;
        RECT 79.565 22.245 79.895 22.615 ;
        RECT 61.085 22.245 61.415 22.615 ;
      LAYER met1 ;
        RECT 170.15 22.28 170.47 22.54 ;
        RECT 133.365 22.295 133.655 22.525 ;
        RECT 131.51 22.34 133.655 22.48 ;
        RECT 131.51 22.28 131.83 22.54 ;
        RECT 79.545 22.295 79.835 22.525 ;
        RECT 79.07 22.34 79.835 22.48 ;
        RECT 79.07 22.28 79.39 22.54 ;
        RECT 61.22 22.68 79.3 22.82 ;
        RECT 79.16 22.28 79.3 22.82 ;
        RECT 61.145 22.295 61.435 22.525 ;
        RECT 61.22 22.295 61.36 22.82 ;
      LAYER met4 ;
        RECT 170.835 22.205 171.165 22.535 ;
        RECT 170.835 0.855 171.165 1.185 ;
        RECT 170.85 0.855 171.15 22.535 ;
      LAYER met3 ;
        RECT 189.465 0.855 189.795 1.185 ;
        RECT 170.81 0.87 189.795 1.17 ;
        RECT 170.81 0.86 171.19 1.18 ;
        RECT 170.81 22.21 171.19 22.53 ;
        RECT 79.065 22.22 171.19 22.52 ;
        RECT 170.145 22.205 170.475 22.535 ;
        RECT 131.505 22.205 131.835 22.535 ;
        RECT 79.065 22.205 79.395 22.535 ;
      LAYER met2 ;
        RECT 189.49 0.835 189.77 1.205 ;
        RECT 189.56 0 189.7 1.205 ;
        RECT 170.17 22.185 170.45 22.555 ;
        RECT 170.18 22.185 170.44 22.57 ;
        RECT 131.53 22.185 131.81 22.555 ;
        RECT 131.54 22.185 131.8 22.57 ;
        RECT 79.09 22.185 79.37 22.555 ;
        RECT 79.1 22.185 79.36 22.57 ;
      LAYER via3 ;
        RECT 170.9 22.27 171.1 22.47 ;
        RECT 170.9 0.92 171.1 1.12 ;
      LAYER via ;
        RECT 79.155 22.335 79.305 22.485 ;
        RECT 131.595 22.335 131.745 22.485 ;
        RECT 170.235 22.335 170.385 22.485 ;
      LAYER mcon ;
        RECT 61.205 22.325 61.375 22.495 ;
        RECT 79.605 22.325 79.775 22.495 ;
        RECT 133.425 22.325 133.595 22.495 ;
        RECT 170.225 22.325 170.395 22.495 ;
      LAYER via2 ;
        RECT 79.13 22.27 79.33 22.47 ;
        RECT 131.57 22.27 131.77 22.47 ;
        RECT 170.21 22.27 170.41 22.47 ;
        RECT 189.53 0.92 189.73 1.12 ;
    END
  END clk
  PIN comp_in
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 171.885 22.275 172.245 22.855 ;
        RECT 170.405 13.795 170.85 13.995 ;
        RECT 119.965 33.155 120.295 33.405 ;
      LAYER met1 ;
        RECT 172.005 22.635 172.295 22.865 ;
        RECT 170.24 22.68 172.295 22.82 ;
        RECT 170.15 22.96 170.47 23.22 ;
        RECT 170.24 22.68 170.38 23.22 ;
        RECT 170.15 13.795 170.685 14.025 ;
        RECT 170.15 13.78 170.47 14.04 ;
        RECT 170.15 32.82 170.47 33.08 ;
        RECT 120.025 33.22 170.38 33.36 ;
        RECT 170.24 32.82 170.38 33.36 ;
        RECT 120.025 33.175 120.315 33.405 ;
      LAYER met2 ;
        RECT 170.24 9.42 170.84 9.56 ;
        RECT 170.7 0 170.84 9.56 ;
        RECT 170.18 32.79 170.44 33.11 ;
        RECT 170.18 22.93 170.44 23.25 ;
        RECT 170.18 13.75 170.44 14.07 ;
        RECT 170.24 22.93 170.38 33.11 ;
        RECT 169.78 16.56 170.38 16.7 ;
        RECT 170.24 9.42 170.38 16.7 ;
        RECT 169.78 23.02 170.44 23.16 ;
        RECT 169.78 16.56 169.92 23.16 ;
      LAYER via ;
        RECT 170.235 32.875 170.385 33.025 ;
        RECT 170.235 23.015 170.385 23.165 ;
        RECT 170.235 13.835 170.385 13.985 ;
      LAYER mcon ;
        RECT 120.085 33.205 120.255 33.375 ;
        RECT 170.455 13.825 170.625 13.995 ;
        RECT 172.065 22.665 172.235 22.835 ;
    END
  END comp_in
  PIN out[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.575 15.695 23.745 17.905 ;
        RECT 21.055 17.255 23.745 17.425 ;
        RECT 23.49 16.545 23.745 17.425 ;
        RECT 21.055 16.545 23.745 16.715 ;
        RECT 22.735 17.255 22.905 17.905 ;
        RECT 22.735 15.695 22.905 16.715 ;
        RECT 21.895 17.255 22.065 17.905 ;
        RECT 21.895 15.695 22.065 16.715 ;
        RECT 21.055 17.255 21.225 17.905 ;
        RECT 21.055 15.695 21.225 16.715 ;
      LAYER met1 ;
        RECT 21.125 16.515 21.415 16.745 ;
        RECT 10.07 16.56 21.415 16.7 ;
        RECT 10.07 16.5 10.39 16.76 ;
      LAYER met2 ;
        RECT 10.1 16.47 10.36 16.79 ;
        RECT 10.16 15.54 10.3 16.79 ;
        RECT 9.7 9.42 10.3 9.56 ;
        RECT 10.16 0 10.3 9.56 ;
        RECT 9.7 15.54 10.3 15.68 ;
        RECT 9.7 9.42 9.84 15.68 ;
      LAYER via ;
        RECT 10.155 16.555 10.305 16.705 ;
      LAYER mcon ;
        RECT 21.185 16.545 21.355 16.715 ;
    END
  END out[15]
  PIN out[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 25.415 23.855 25.585 26.065 ;
        RECT 22.895 25.045 25.585 25.215 ;
        RECT 25.33 24.335 25.585 25.215 ;
        RECT 22.895 24.335 25.585 24.505 ;
        RECT 24.575 25.045 24.745 26.065 ;
        RECT 24.575 23.855 24.745 24.505 ;
        RECT 23.735 25.045 23.905 26.065 ;
        RECT 23.735 23.855 23.905 24.505 ;
        RECT 22.895 25.045 23.065 26.065 ;
        RECT 22.895 23.855 23.065 24.505 ;
      LAYER met1 ;
        RECT 22.965 25.015 23.255 25.245 ;
        RECT 18.35 25.06 23.255 25.2 ;
        RECT 18.35 25 18.67 25.26 ;
      LAYER met2 ;
        RECT 19.82 0 19.96 0.485 ;
        RECT 18.44 0.34 19.96 0.48 ;
        RECT 18.38 24.97 18.64 25.29 ;
        RECT 18.44 0.34 18.58 25.29 ;
      LAYER via ;
        RECT 18.435 25.055 18.585 25.205 ;
      LAYER mcon ;
        RECT 23.025 25.045 23.195 25.215 ;
    END
  END out[16]
  PIN out[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 34.155 15.695 34.325 17.905 ;
        RECT 31.635 17.255 34.325 17.425 ;
        RECT 34.07 16.545 34.325 17.425 ;
        RECT 31.635 16.545 34.325 16.715 ;
        RECT 33.315 17.255 33.485 17.905 ;
        RECT 33.315 15.695 33.485 16.715 ;
        RECT 32.475 17.255 32.645 17.905 ;
        RECT 32.475 15.695 32.645 16.715 ;
        RECT 31.635 17.255 31.805 17.905 ;
        RECT 31.635 15.695 31.805 16.715 ;
      LAYER met1 ;
        RECT 31.705 16.515 31.995 16.745 ;
        RECT 29.39 16.56 31.995 16.7 ;
        RECT 29.39 16.5 29.71 16.76 ;
      LAYER met2 ;
        RECT 29.42 16.47 29.68 16.79 ;
        RECT 29.48 0 29.62 16.79 ;
      LAYER via ;
        RECT 29.475 16.555 29.625 16.705 ;
      LAYER mcon ;
        RECT 31.765 16.545 31.935 16.715 ;
    END
  END out[17]
  PIN out[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 38.795 28.135 38.965 28.785 ;
        RECT 36.275 27.425 38.965 27.595 ;
        RECT 38.795 26.575 38.965 27.595 ;
        RECT 36.275 28.135 38.965 28.305 ;
        RECT 37.955 28.135 38.125 28.785 ;
        RECT 37.955 26.575 38.125 27.595 ;
        RECT 37.115 28.135 37.285 28.785 ;
        RECT 37.115 26.575 37.285 27.595 ;
        RECT 36.275 27.425 36.53 28.305 ;
        RECT 36.275 26.575 36.445 28.785 ;
      LAYER met1 ;
        RECT 37.67 27.38 37.99 27.64 ;
      LAYER met2 ;
        RECT 37.76 9.08 38.82 9.22 ;
        RECT 38.68 0 38.82 9.22 ;
        RECT 37.7 27.35 37.96 27.67 ;
        RECT 37.76 9.08 37.9 27.67 ;
      LAYER via ;
        RECT 37.755 27.435 37.905 27.585 ;
      LAYER mcon ;
        RECT 37.745 27.425 37.915 27.595 ;
    END
  END out[18]
  PIN out[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 39.255 17.255 39.425 17.905 ;
        RECT 36.735 16.545 39.425 16.715 ;
        RECT 39.255 15.695 39.425 16.715 ;
        RECT 36.735 17.255 39.425 17.425 ;
        RECT 38.415 17.255 38.585 17.905 ;
        RECT 38.415 15.695 38.585 16.715 ;
        RECT 37.575 17.255 37.745 17.905 ;
        RECT 37.575 15.695 37.745 16.715 ;
        RECT 36.735 16.545 36.99 17.425 ;
        RECT 36.735 15.695 36.905 17.905 ;
      LAYER met1 ;
        RECT 48.25 0.52 48.57 0.78 ;
        RECT 40.43 0.58 48.57 0.72 ;
        RECT 40.43 0.52 40.75 0.78 ;
        RECT 40.43 16.16 40.75 16.42 ;
        RECT 39.065 16.56 40.66 16.7 ;
        RECT 40.52 16.16 40.66 16.7 ;
        RECT 39.065 16.515 39.355 16.745 ;
      LAYER met2 ;
        RECT 48.28 0.49 48.54 0.81 ;
        RECT 48.34 0 48.48 0.81 ;
        RECT 40.46 16.13 40.72 16.45 ;
        RECT 40.46 0.49 40.72 0.81 ;
        RECT 40.52 0.49 40.66 16.45 ;
      LAYER via ;
        RECT 40.515 16.215 40.665 16.365 ;
        RECT 40.515 0.575 40.665 0.725 ;
        RECT 48.335 0.575 48.485 0.725 ;
      LAYER mcon ;
        RECT 39.125 16.545 39.295 16.715 ;
    END
  END out[19]
  PIN out[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 70.035 23.855 70.205 26.065 ;
        RECT 67.515 25.045 70.205 25.215 ;
        RECT 69.95 24.335 70.205 25.215 ;
        RECT 69.945 24.335 70.205 24.535 ;
        RECT 67.515 24.335 70.205 24.505 ;
        RECT 69.195 25.045 69.365 26.065 ;
        RECT 69.195 23.855 69.365 24.505 ;
        RECT 68.355 25.045 68.525 26.065 ;
        RECT 68.355 23.855 68.525 24.505 ;
        RECT 67.515 25.045 67.685 26.065 ;
        RECT 67.515 23.855 67.685 24.505 ;
      LAYER met1 ;
        RECT 69.885 24.335 70.175 24.565 ;
        RECT 67.66 24.38 70.175 24.52 ;
        RECT 67.66 24.04 67.8 24.52 ;
        RECT 64.44 24.04 67.8 24.18 ;
        RECT 58 24.21 64.58 24.35 ;
        RECT 64.44 24.04 64.58 24.35 ;
        RECT 58 24.04 58.14 24.35 ;
        RECT 56.99 24.04 58.14 24.18 ;
        RECT 56.99 23.98 57.31 24.24 ;
      LAYER met2 ;
        RECT 57.02 24.04 57.68 24.18 ;
        RECT 57.54 12.82 57.68 24.18 ;
        RECT 57.08 9.42 57.68 9.56 ;
        RECT 57.54 0 57.68 9.56 ;
        RECT 57.08 12.82 57.68 12.96 ;
        RECT 57.02 23.95 57.28 24.27 ;
        RECT 57.08 9.42 57.22 12.96 ;
      LAYER via ;
        RECT 57.075 24.035 57.225 24.185 ;
      LAYER mcon ;
        RECT 69.945 24.365 70.115 24.535 ;
    END
  END out[20]
  PIN out[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 70.035 12.975 70.205 15.185 ;
        RECT 67.515 14.165 70.205 14.335 ;
        RECT 69.95 13.455 70.205 14.335 ;
        RECT 67.515 13.455 70.205 13.625 ;
        RECT 69.195 14.165 69.365 15.185 ;
        RECT 69.195 12.975 69.365 13.625 ;
        RECT 68.355 14.165 68.525 15.185 ;
        RECT 68.355 12.975 68.525 13.625 ;
        RECT 67.515 14.165 67.685 15.185 ;
        RECT 67.515 12.975 67.685 13.625 ;
      LAYER met1 ;
        RECT 68.03 14.12 68.35 14.38 ;
      LAYER met2 ;
        RECT 68.06 14.09 68.32 14.41 ;
        RECT 68.12 2.28 68.26 14.41 ;
        RECT 67.2 2.28 68.26 2.42 ;
        RECT 67.2 0 67.34 2.42 ;
      LAYER via ;
        RECT 68.115 14.175 68.265 14.325 ;
      LAYER mcon ;
        RECT 68.105 14.165 68.275 14.335 ;
    END
  END out[21]
  PIN out[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 78.315 10.255 78.485 12.465 ;
        RECT 75.795 11.815 78.485 11.985 ;
        RECT 78.23 11.105 78.485 11.985 ;
        RECT 75.795 11.105 78.485 11.275 ;
        RECT 77.475 11.815 77.645 12.465 ;
        RECT 77.475 10.255 77.645 11.275 ;
        RECT 76.635 11.815 76.805 12.465 ;
        RECT 76.635 10.255 76.805 11.275 ;
        RECT 75.795 11.815 75.965 12.465 ;
        RECT 75.795 10.255 75.965 11.275 ;
      LAYER met1 ;
        RECT 79.07 11.06 79.39 11.32 ;
        RECT 78.165 11.12 79.39 11.26 ;
        RECT 78.165 11.075 78.455 11.305 ;
      LAYER met2 ;
        RECT 79.1 11.03 79.36 11.35 ;
        RECT 79.16 9.08 79.3 11.35 ;
        RECT 77.78 9.08 79.3 9.22 ;
        RECT 77.78 0.34 77.92 9.22 ;
        RECT 76.4 0.34 77.92 0.48 ;
        RECT 76.4 0 76.54 0.485 ;
      LAYER via ;
        RECT 79.155 11.115 79.305 11.265 ;
      LAYER mcon ;
        RECT 78.225 11.105 78.395 11.275 ;
    END
  END out[22]
  PIN out[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 95.795 10.255 95.965 12.465 ;
        RECT 93.275 11.815 95.965 11.985 ;
        RECT 95.71 11.105 95.965 11.985 ;
        RECT 93.275 11.105 95.965 11.275 ;
        RECT 94.955 11.815 95.125 12.465 ;
        RECT 94.955 10.255 95.125 11.275 ;
        RECT 94.115 11.815 94.285 12.465 ;
        RECT 94.115 10.255 94.285 11.275 ;
        RECT 93.275 11.815 93.445 12.465 ;
        RECT 93.275 10.255 93.445 11.275 ;
      LAYER met1 ;
        RECT 93.345 11.075 93.635 11.305 ;
        RECT 92.87 11.12 93.635 11.26 ;
        RECT 92.87 11.06 93.19 11.32 ;
        RECT 92.87 0.52 93.19 0.78 ;
        RECT 85.97 0.58 93.19 0.72 ;
        RECT 85.97 0.52 86.29 0.78 ;
      LAYER met2 ;
        RECT 92.9 11.03 93.16 11.35 ;
        RECT 92.9 0.49 93.16 0.81 ;
        RECT 92.96 0.49 93.1 11.35 ;
        RECT 86 0.49 86.26 0.81 ;
        RECT 86.06 0 86.2 0.81 ;
      LAYER via ;
        RECT 86.055 0.575 86.205 0.725 ;
        RECT 92.955 11.115 93.105 11.265 ;
        RECT 92.955 0.575 93.105 0.725 ;
      LAYER mcon ;
        RECT 93.405 11.105 93.575 11.275 ;
    END
  END out[23]
  PIN out[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 101.775 10.255 101.945 12.465 ;
        RECT 99.255 11.815 101.945 11.985 ;
        RECT 101.69 11.105 101.945 11.985 ;
        RECT 99.255 11.105 101.945 11.275 ;
        RECT 100.935 11.815 101.105 12.465 ;
        RECT 100.935 10.255 101.105 11.275 ;
        RECT 100.095 11.815 100.265 12.465 ;
        RECT 100.095 10.255 100.265 11.275 ;
        RECT 99.255 11.815 99.425 12.465 ;
        RECT 99.255 10.255 99.425 11.275 ;
      LAYER met1 ;
        RECT 99.325 11.075 99.615 11.305 ;
        RECT 95.63 11.12 99.615 11.26 ;
        RECT 95.63 11.06 95.95 11.32 ;
      LAYER met2 ;
        RECT 95.66 11.03 95.92 11.35 ;
        RECT 95.26 11.12 95.92 11.26 ;
        RECT 95.26 0 95.4 11.26 ;
      LAYER via ;
        RECT 95.715 11.115 95.865 11.265 ;
      LAYER mcon ;
        RECT 99.385 11.105 99.555 11.275 ;
    END
  END out[24]
  PIN out[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 107.755 12.975 107.925 15.185 ;
        RECT 105.235 14.165 107.925 14.335 ;
        RECT 107.67 13.455 107.925 14.335 ;
        RECT 105.235 13.455 107.925 13.625 ;
        RECT 106.915 14.165 107.085 15.185 ;
        RECT 106.915 12.975 107.085 13.625 ;
        RECT 106.075 14.165 106.245 15.185 ;
        RECT 106.075 12.975 106.245 13.625 ;
        RECT 105.235 14.165 105.405 15.185 ;
        RECT 105.235 12.975 105.405 13.625 ;
      LAYER met1 ;
        RECT 105.305 14.135 105.595 14.365 ;
        RECT 103.91 14.18 105.595 14.32 ;
        RECT 103.91 14.12 104.23 14.38 ;
      LAYER met2 ;
        RECT 104.92 0 105.06 0.485 ;
        RECT 104 0.34 105.06 0.48 ;
        RECT 103.94 14.09 104.2 14.41 ;
        RECT 104 0.34 104.14 14.41 ;
      LAYER via ;
        RECT 103.995 14.175 104.145 14.325 ;
      LAYER mcon ;
        RECT 105.365 14.165 105.535 14.335 ;
    END
  END out[25]
  PIN out[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 113.775 14.165 113.945 15.185 ;
        RECT 111.255 13.455 113.945 13.625 ;
        RECT 113.775 12.975 113.945 13.625 ;
        RECT 111.255 14.165 113.945 14.335 ;
        RECT 112.935 14.165 113.105 15.185 ;
        RECT 112.935 12.975 113.105 13.625 ;
        RECT 112.095 14.165 112.265 15.185 ;
        RECT 112.095 12.975 112.265 13.625 ;
        RECT 111.255 13.455 111.51 14.335 ;
        RECT 111.255 12.975 111.425 15.185 ;
      LAYER met1 ;
        RECT 114.95 14.12 115.27 14.38 ;
        RECT 113.585 14.18 115.27 14.32 ;
        RECT 113.585 14.135 113.875 14.365 ;
      LAYER met2 ;
        RECT 114.98 14.09 115.24 14.41 ;
        RECT 115.04 9.08 115.18 14.41 ;
        RECT 114.12 9.08 115.18 9.22 ;
        RECT 114.12 0 114.26 9.22 ;
      LAYER via ;
        RECT 115.035 14.175 115.185 14.325 ;
      LAYER mcon ;
        RECT 113.645 14.165 113.815 14.335 ;
    END
  END out[26]
  PIN out[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 121.595 11.815 121.765 12.465 ;
        RECT 119.075 11.105 121.765 11.275 ;
        RECT 121.595 10.255 121.765 11.275 ;
        RECT 119.075 11.815 121.765 11.985 ;
        RECT 120.755 11.815 120.925 12.465 ;
        RECT 120.755 10.255 120.925 11.275 ;
        RECT 119.915 11.815 120.085 12.465 ;
        RECT 119.915 10.255 120.085 11.275 ;
        RECT 119.075 11.105 119.33 11.985 ;
        RECT 119.075 10.255 119.245 12.465 ;
      LAYER met1 ;
        RECT 123.23 11.06 123.55 11.32 ;
        RECT 121.405 11.12 123.55 11.26 ;
        RECT 121.405 11.075 121.695 11.305 ;
      LAYER met2 ;
        RECT 123.32 9.08 123.92 9.22 ;
        RECT 123.78 0 123.92 9.22 ;
        RECT 123.26 11.03 123.52 11.35 ;
        RECT 123.32 9.08 123.46 11.35 ;
      LAYER via ;
        RECT 123.315 11.115 123.465 11.265 ;
      LAYER mcon ;
        RECT 121.465 11.105 121.635 11.275 ;
    END
  END out[27]
  PIN out[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 137.195 12.975 137.365 15.185 ;
        RECT 134.675 14.165 137.365 14.335 ;
        RECT 137.11 13.455 137.365 14.335 ;
        RECT 134.675 13.455 137.365 13.625 ;
        RECT 136.355 14.165 136.525 15.185 ;
        RECT 136.355 12.975 136.525 13.625 ;
        RECT 135.515 14.165 135.685 15.185 ;
        RECT 135.515 12.975 135.685 13.625 ;
        RECT 134.675 14.165 134.845 15.185 ;
        RECT 134.675 12.975 134.845 13.625 ;
      LAYER met1 ;
        RECT 134.745 14.135 135.035 14.365 ;
        RECT 134.27 14.18 135.035 14.32 ;
        RECT 134.27 14.12 134.59 14.38 ;
      LAYER met2 ;
        RECT 134.3 14.09 134.56 14.41 ;
        RECT 134.36 0.34 134.5 14.41 ;
        RECT 132.98 0.34 134.5 0.48 ;
        RECT 132.98 0 133.12 0.485 ;
      LAYER via ;
        RECT 134.355 14.175 134.505 14.325 ;
      LAYER mcon ;
        RECT 134.805 14.165 134.975 14.335 ;
    END
  END out[28]
  PIN out[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 142.755 14.165 142.925 15.185 ;
        RECT 140.235 13.455 142.925 13.625 ;
        RECT 142.755 12.975 142.925 13.625 ;
        RECT 140.235 14.165 142.925 14.335 ;
        RECT 141.915 14.165 142.085 15.185 ;
        RECT 141.915 12.975 142.085 13.625 ;
        RECT 141.075 14.165 141.245 15.185 ;
        RECT 141.075 12.975 141.245 13.625 ;
        RECT 140.235 13.455 140.49 14.335 ;
        RECT 140.235 12.975 140.405 15.185 ;
      LAYER met1 ;
        RECT 142.55 14.12 142.87 14.38 ;
      LAYER met2 ;
        RECT 142.58 14.09 142.84 14.41 ;
        RECT 142.64 0 142.78 14.41 ;
      LAYER via ;
        RECT 142.635 14.175 142.785 14.325 ;
      LAYER mcon ;
        RECT 142.625 14.165 142.795 14.335 ;
    END
  END out[29]
  PIN out[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 152.835 10.255 153.005 12.465 ;
        RECT 150.315 11.815 153.005 11.985 ;
        RECT 152.75 11.105 153.005 11.985 ;
        RECT 150.315 11.105 153.005 11.275 ;
        RECT 151.995 11.815 152.165 12.465 ;
        RECT 151.995 10.255 152.165 11.275 ;
        RECT 151.155 11.815 151.325 12.465 ;
        RECT 151.155 10.255 151.325 11.275 ;
        RECT 150.315 11.815 150.485 12.465 ;
        RECT 150.315 10.255 150.485 11.275 ;
      LAYER met1 ;
        RECT 153.59 11.06 153.91 11.32 ;
        RECT 152.685 11.12 153.91 11.26 ;
        RECT 152.685 11.075 152.975 11.305 ;
      LAYER met2 ;
        RECT 153.62 11.03 153.88 11.35 ;
        RECT 153.68 0.92 153.82 11.35 ;
        RECT 151.84 0.92 153.82 1.06 ;
        RECT 151.84 0 151.98 1.06 ;
      LAYER via ;
        RECT 153.675 11.115 153.825 11.265 ;
      LAYER mcon ;
        RECT 152.745 11.105 152.915 11.275 ;
    END
  END out[30]
  PIN out[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 167.555 10.255 167.725 12.465 ;
        RECT 165.035 11.815 167.725 11.985 ;
        RECT 167.47 11.105 167.725 11.985 ;
        RECT 165.035 11.105 167.725 11.275 ;
        RECT 166.715 11.815 166.885 12.465 ;
        RECT 166.715 10.255 166.885 11.275 ;
        RECT 165.875 11.815 166.045 12.465 ;
        RECT 165.875 10.255 166.045 11.275 ;
        RECT 165.035 11.815 165.205 12.465 ;
        RECT 165.035 10.255 165.205 11.275 ;
      LAYER met1 ;
        RECT 165.105 11.075 165.395 11.305 ;
        RECT 161.87 11.12 165.395 11.26 ;
        RECT 161.87 11.06 162.19 11.32 ;
      LAYER met2 ;
        RECT 161.9 11.03 162.16 11.35 ;
        RECT 161.96 9.76 162.1 11.35 ;
        RECT 161.5 9.76 162.1 9.9 ;
        RECT 161.5 0 161.64 9.9 ;
      LAYER via ;
        RECT 161.955 11.115 162.105 11.265 ;
      LAYER mcon ;
        RECT 165.165 11.105 165.335 11.275 ;
    END
  END out[31]
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 173.265 18.905 173.625 19.485 ;
        RECT 171.02 13.795 171.37 14.005 ;
      LAYER met1 ;
        RECT 180.27 9.36 180.59 9.62 ;
        RECT 179.44 9.42 180.59 9.56 ;
        RECT 179.44 8.74 179.58 9.56 ;
        RECT 174.38 8.74 179.58 8.88 ;
        RECT 173.37 9.42 174.52 9.56 ;
        RECT 174.38 8.74 174.52 9.56 ;
        RECT 173.37 9.36 173.69 9.62 ;
        RECT 173.385 19.235 173.675 19.465 ;
        RECT 172.91 19.28 173.675 19.42 ;
        RECT 172.91 19.22 173.23 19.48 ;
        RECT 172.91 13.78 173.23 14.04 ;
        RECT 171.085 13.84 173.23 13.98 ;
        RECT 171.085 13.795 171.375 14.025 ;
      LAYER met2 ;
        RECT 180.3 9.33 180.56 9.65 ;
        RECT 180.36 0 180.5 9.65 ;
        RECT 173.4 9.33 173.66 9.65 ;
        RECT 172.94 19.28 173.6 19.42 ;
        RECT 173.46 9.33 173.6 19.42 ;
        RECT 172.94 13.84 173.6 13.98 ;
        RECT 172.94 19.19 173.2 19.51 ;
        RECT 172.94 13.75 173.2 14.07 ;
      LAYER via ;
        RECT 172.995 19.275 173.145 19.425 ;
        RECT 172.995 13.835 173.145 13.985 ;
        RECT 173.455 9.415 173.605 9.565 ;
        RECT 180.355 9.415 180.505 9.565 ;
      LAYER mcon ;
        RECT 171.145 13.825 171.315 13.995 ;
        RECT 173.445 19.265 173.615 19.435 ;
    END
  END rst
  PIN out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 23.575 12.975 23.745 15.185 ;
        RECT 21.055 14.165 23.745 14.335 ;
        RECT 23.49 13.455 23.745 14.335 ;
        RECT 21.055 13.455 23.745 13.625 ;
        RECT 22.735 14.165 22.905 15.185 ;
        RECT 22.735 12.975 22.905 13.625 ;
        RECT 21.895 14.165 22.065 15.185 ;
        RECT 21.895 12.975 22.065 13.625 ;
        RECT 21.055 14.165 21.225 15.185 ;
        RECT 21.055 12.975 21.225 13.625 ;
      LAYER met1 ;
        RECT 21.125 14.135 21.415 14.365 ;
        RECT 15.59 14.18 21.415 14.32 ;
        RECT 15.59 14.12 15.91 14.38 ;
      LAYER met4 ;
        RECT 10.065 1.465 10.395 1.795 ;
        RECT 10.08 0 10.38 1.795 ;
      LAYER met3 ;
        RECT 15.585 1.465 15.915 1.795 ;
        RECT 10.04 1.48 15.915 1.78 ;
        RECT 10.04 1.47 10.42 1.79 ;
      LAYER met2 ;
        RECT 15.61 1.445 15.89 1.815 ;
        RECT 15.62 14.09 15.88 14.41 ;
        RECT 15.68 1.445 15.82 14.41 ;
      LAYER via3 ;
        RECT 10.13 1.53 10.33 1.73 ;
      LAYER via ;
        RECT 15.675 14.175 15.825 14.325 ;
      LAYER mcon ;
        RECT 21.185 14.165 21.355 14.335 ;
      LAYER via2 ;
        RECT 15.65 1.53 15.85 1.73 ;
    END
  END out[0]
  PIN out[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 142.715 10.255 142.885 12.465 ;
        RECT 140.195 11.815 142.885 11.985 ;
        RECT 142.63 11.105 142.885 11.985 ;
        RECT 140.195 11.105 142.885 11.275 ;
        RECT 141.875 11.815 142.045 12.465 ;
        RECT 141.875 10.255 142.045 11.275 ;
        RECT 141.035 11.815 141.205 12.465 ;
        RECT 141.035 10.255 141.205 11.275 ;
        RECT 140.195 11.815 140.365 12.465 ;
        RECT 140.195 10.255 140.365 11.275 ;
      LAYER met1 ;
        RECT 140.265 11.075 140.555 11.305 ;
        RECT 137.03 11.12 140.555 11.26 ;
        RECT 137.03 11.06 137.35 11.32 ;
      LAYER met4 ;
        RECT 138.405 0.855 138.735 1.185 ;
        RECT 138.42 0 138.72 1.185 ;
      LAYER met3 ;
        RECT 138.38 0.86 138.76 1.18 ;
        RECT 137.025 0.87 138.76 1.17 ;
        RECT 137.025 0.855 137.355 1.185 ;
      LAYER met2 ;
        RECT 137.05 0.835 137.33 1.205 ;
        RECT 137.06 11.03 137.32 11.35 ;
        RECT 137.12 0.835 137.26 11.35 ;
      LAYER via3 ;
        RECT 138.47 0.92 138.67 1.12 ;
      LAYER via ;
        RECT 137.115 11.115 137.265 11.265 ;
      LAYER mcon ;
        RECT 140.325 11.105 140.495 11.275 ;
      LAYER via2 ;
        RECT 137.09 0.92 137.29 1.12 ;
    END
  END out[10]
  PIN out[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 151.035 25.045 151.205 26.065 ;
        RECT 148.515 24.335 151.205 24.505 ;
        RECT 151.035 23.855 151.205 24.505 ;
        RECT 148.515 25.045 151.205 25.215 ;
        RECT 150.195 25.045 150.365 26.065 ;
        RECT 150.195 23.855 150.365 24.505 ;
        RECT 149.355 25.045 149.525 26.065 ;
        RECT 149.355 23.855 149.525 24.505 ;
        RECT 148.515 24.335 148.77 25.215 ;
        RECT 148.515 23.855 148.685 26.065 ;
      LAYER met1 ;
        RECT 150.83 25 151.15 25.26 ;
      LAYER met4 ;
        RECT 151.515 8.785 151.845 9.115 ;
        RECT 151.53 0 151.83 9.115 ;
      LAYER met3 ;
        RECT 151.285 8.79 151.87 9.11 ;
        RECT 151.285 8.785 151.615 9.115 ;
        RECT 151.07 8.8 151.87 9.1 ;
      LAYER met2 ;
        RECT 151.31 8.765 151.59 9.135 ;
        RECT 150.92 17.24 151.52 17.38 ;
        RECT 151.38 8.765 151.52 17.38 ;
        RECT 150.86 24.97 151.12 25.29 ;
        RECT 150.92 17.24 151.06 25.29 ;
      LAYER via3 ;
        RECT 151.58 8.85 151.78 9.05 ;
      LAYER via ;
        RECT 150.915 25.055 151.065 25.205 ;
      LAYER mcon ;
        RECT 150.905 25.045 151.075 25.215 ;
      LAYER via2 ;
        RECT 151.35 8.85 151.55 9.05 ;
    END
  END out[11]
  PIN out[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 166.635 15.695 166.805 17.905 ;
        RECT 164.115 17.255 166.805 17.425 ;
        RECT 166.55 16.545 166.805 17.425 ;
        RECT 164.115 16.545 166.805 16.715 ;
        RECT 165.795 17.255 165.965 17.905 ;
        RECT 165.795 15.695 165.965 16.715 ;
        RECT 164.955 17.255 165.125 17.905 ;
        RECT 164.955 15.695 165.125 16.715 ;
        RECT 164.115 17.255 164.285 17.905 ;
        RECT 164.115 15.695 164.285 16.715 ;
      LAYER met1 ;
        RECT 164.63 16.5 164.95 16.76 ;
      LAYER met4 ;
        RECT 163.935 3.295 164.265 3.625 ;
        RECT 163.95 0 164.25 3.625 ;
      LAYER met3 ;
        RECT 164.625 3.295 164.955 3.625 ;
        RECT 163.91 3.31 164.955 3.61 ;
        RECT 163.91 3.3 164.29 3.62 ;
      LAYER met2 ;
        RECT 164.65 3.275 164.93 3.645 ;
        RECT 164.66 16.47 164.92 16.79 ;
        RECT 164.72 3.275 164.86 16.79 ;
      LAYER via3 ;
        RECT 164 3.36 164.2 3.56 ;
      LAYER via ;
        RECT 164.715 16.555 164.865 16.705 ;
      LAYER mcon ;
        RECT 164.705 16.545 164.875 16.715 ;
      LAYER via2 ;
        RECT 164.69 3.36 164.89 3.56 ;
    END
  END out[12]
  PIN out[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 181.355 15.695 181.525 17.905 ;
        RECT 178.835 17.255 181.525 17.425 ;
        RECT 181.27 16.545 181.525 17.425 ;
        RECT 178.835 16.545 181.525 16.715 ;
        RECT 180.515 17.255 180.685 17.905 ;
        RECT 180.515 15.695 180.685 16.715 ;
        RECT 179.675 17.255 179.845 17.905 ;
        RECT 179.675 15.695 179.845 16.715 ;
        RECT 178.835 17.255 179.005 17.905 ;
        RECT 178.835 15.695 179.005 16.715 ;
      LAYER met1 ;
        RECT 178.905 16.515 179.195 16.745 ;
        RECT 178.43 16.56 179.195 16.7 ;
        RECT 178.43 16.5 178.75 16.76 ;
      LAYER met4 ;
        RECT 177.045 3.905 177.375 4.235 ;
        RECT 177.06 0 177.36 4.235 ;
      LAYER met3 ;
        RECT 178.425 3.905 178.755 4.235 ;
        RECT 177.02 3.92 178.755 4.22 ;
        RECT 177.02 3.91 177.4 4.23 ;
      LAYER met2 ;
        RECT 178.45 3.885 178.73 4.255 ;
        RECT 178.46 16.47 178.72 16.79 ;
        RECT 178.52 3.885 178.66 16.79 ;
      LAYER via3 ;
        RECT 177.11 3.97 177.31 4.17 ;
      LAYER via ;
        RECT 178.515 16.555 178.665 16.705 ;
      LAYER mcon ;
        RECT 178.965 16.545 179.135 16.715 ;
      LAYER via2 ;
        RECT 178.49 3.97 178.69 4.17 ;
    END
  END out[13]
  PIN out[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 184.575 23.855 184.745 26.065 ;
        RECT 182.055 25.045 184.745 25.215 ;
        RECT 184.49 24.335 184.745 25.215 ;
        RECT 184.485 24.335 184.745 24.535 ;
        RECT 182.055 24.335 184.745 24.505 ;
        RECT 183.735 25.045 183.905 26.065 ;
        RECT 183.735 23.855 183.905 24.505 ;
        RECT 182.895 25.045 183.065 26.065 ;
        RECT 182.895 23.855 183.065 24.505 ;
        RECT 182.055 25.045 182.225 26.065 ;
        RECT 182.055 23.855 182.225 24.505 ;
      LAYER met1 ;
        RECT 186.71 24.32 187.03 24.58 ;
        RECT 184.425 24.38 187.03 24.52 ;
        RECT 184.425 24.335 184.715 24.565 ;
      LAYER met4 ;
        RECT 189.465 5.125 189.795 5.455 ;
        RECT 189.48 0 189.78 5.455 ;
      LAYER met3 ;
        RECT 189.44 5.13 189.82 5.45 ;
        RECT 186.705 5.14 189.82 5.44 ;
        RECT 186.705 5.125 187.035 5.455 ;
      LAYER met2 ;
        RECT 186.73 5.105 187.01 5.475 ;
        RECT 186.74 24.29 187 24.61 ;
        RECT 186.8 5.105 186.94 24.61 ;
      LAYER via3 ;
        RECT 189.53 5.19 189.73 5.39 ;
      LAYER via ;
        RECT 186.795 24.375 186.945 24.525 ;
      LAYER mcon ;
        RECT 184.485 24.365 184.655 24.535 ;
      LAYER via2 ;
        RECT 186.77 5.19 186.97 5.39 ;
    END
  END out[14]
  PIN out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 34.155 10.255 34.325 12.465 ;
        RECT 31.635 11.815 34.325 11.985 ;
        RECT 34.07 11.105 34.325 11.985 ;
        RECT 31.635 11.105 34.325 11.275 ;
        RECT 33.315 11.815 33.485 12.465 ;
        RECT 33.315 10.255 33.485 11.275 ;
        RECT 32.475 11.815 32.645 12.465 ;
        RECT 32.475 10.255 32.645 11.275 ;
        RECT 31.635 11.815 31.805 12.465 ;
        RECT 31.635 10.255 31.805 11.275 ;
      LAYER met1 ;
        RECT 31.705 11.075 31.995 11.305 ;
        RECT 26.63 11.12 31.995 11.26 ;
        RECT 26.63 11.06 26.95 11.32 ;
      LAYER met4 ;
        RECT 23.175 0.855 23.505 1.185 ;
        RECT 23.19 0 23.49 1.185 ;
      LAYER met3 ;
        RECT 26.625 0.855 26.955 1.185 ;
        RECT 23.15 0.87 26.955 1.17 ;
        RECT 23.15 0.86 23.53 1.18 ;
      LAYER met2 ;
        RECT 26.65 0.835 26.93 1.205 ;
        RECT 26.66 11.03 26.92 11.35 ;
        RECT 26.72 0.835 26.86 11.35 ;
      LAYER via3 ;
        RECT 23.24 0.92 23.44 1.12 ;
      LAYER via ;
        RECT 26.715 11.115 26.865 11.265 ;
      LAYER mcon ;
        RECT 31.765 11.105 31.935 11.275 ;
      LAYER via2 ;
        RECT 26.69 0.92 26.89 1.12 ;
    END
  END out[1]
  PIN out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 36.035 14.165 36.205 15.185 ;
        RECT 33.515 13.455 36.205 13.625 ;
        RECT 36.035 12.975 36.205 13.625 ;
        RECT 33.515 14.165 36.205 14.335 ;
        RECT 35.195 14.165 35.365 15.185 ;
        RECT 35.195 12.975 35.365 13.625 ;
        RECT 34.355 14.165 34.525 15.185 ;
        RECT 34.355 12.975 34.525 13.625 ;
        RECT 33.515 13.455 33.77 14.335 ;
        RECT 33.515 12.975 33.685 15.185 ;
      LAYER met1 ;
        RECT 34.91 14.12 35.23 14.38 ;
      LAYER met4 ;
        RECT 36.285 0.855 36.615 1.185 ;
        RECT 36.3 0 36.6 1.185 ;
      LAYER met3 ;
        RECT 36.26 0.86 36.64 1.18 ;
        RECT 34.905 0.87 36.64 1.17 ;
        RECT 34.905 0.855 35.235 1.185 ;
      LAYER met2 ;
        RECT 34.93 0.835 35.21 1.205 ;
        RECT 34.94 14.09 35.2 14.41 ;
        RECT 35 0.835 35.14 14.41 ;
      LAYER via3 ;
        RECT 36.35 0.92 36.55 1.12 ;
      LAYER via ;
        RECT 34.995 14.175 35.145 14.325 ;
      LAYER mcon ;
        RECT 34.985 14.165 35.155 14.335 ;
      LAYER via2 ;
        RECT 34.97 0.92 35.17 1.12 ;
    END
  END out[2]
  PIN out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 52.095 10.255 52.265 12.465 ;
        RECT 49.575 11.815 52.265 11.985 ;
        RECT 52.01 11.105 52.265 11.985 ;
        RECT 49.575 11.105 52.265 11.275 ;
        RECT 51.255 11.815 51.425 12.465 ;
        RECT 51.255 10.255 51.425 11.275 ;
        RECT 50.415 11.815 50.585 12.465 ;
        RECT 50.415 10.255 50.585 11.275 ;
        RECT 49.575 11.815 49.745 12.465 ;
        RECT 49.575 10.255 49.745 11.275 ;
      LAYER met1 ;
        RECT 49.57 11.075 49.86 11.305 ;
        RECT 49.645 10.44 49.785 11.305 ;
        RECT 48.71 10.44 49.785 10.58 ;
        RECT 48.71 10.38 49.03 10.64 ;
      LAYER met4 ;
        RECT 48.705 10.005 49.035 10.335 ;
        RECT 48.72 0 49.02 10.335 ;
      LAYER met3 ;
        RECT 48.68 10.01 49.06 10.33 ;
        RECT 48.705 10.005 49.035 10.335 ;
        RECT 48.26 10.02 49.06 10.32 ;
      LAYER met2 ;
        RECT 48.73 9.985 49.01 10.355 ;
        RECT 48.74 9.985 49 10.67 ;
      LAYER via3 ;
        RECT 48.77 10.07 48.97 10.27 ;
      LAYER via ;
        RECT 48.795 10.435 48.945 10.585 ;
      LAYER mcon ;
        RECT 49.63 11.105 49.8 11.275 ;
      LAYER via2 ;
        RECT 48.77 10.07 48.97 10.27 ;
    END
  END out[3]
  PIN out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 66.815 10.255 66.985 12.465 ;
        RECT 64.295 11.815 66.985 11.985 ;
        RECT 66.73 11.105 66.985 11.985 ;
        RECT 64.295 11.105 66.985 11.275 ;
        RECT 65.975 11.815 66.145 12.465 ;
        RECT 65.975 10.255 66.145 11.275 ;
        RECT 65.135 11.815 65.305 12.465 ;
        RECT 65.135 10.255 65.305 11.275 ;
        RECT 64.295 11.815 64.465 12.465 ;
        RECT 64.295 10.255 64.465 11.275 ;
      LAYER met1 ;
        RECT 65.27 11.06 65.59 11.32 ;
      LAYER met4 ;
        RECT 61.815 0.855 62.145 1.185 ;
        RECT 61.83 0 62.13 1.185 ;
      LAYER met3 ;
        RECT 65.265 0.855 65.595 1.185 ;
        RECT 61.79 0.87 65.595 1.17 ;
        RECT 61.79 0.86 62.17 1.18 ;
      LAYER met2 ;
        RECT 65.29 0.835 65.57 1.205 ;
        RECT 65.3 11.03 65.56 11.35 ;
        RECT 65.36 0.835 65.5 11.35 ;
      LAYER via3 ;
        RECT 61.88 0.92 62.08 1.12 ;
      LAYER via ;
        RECT 65.355 11.115 65.505 11.265 ;
      LAYER mcon ;
        RECT 65.345 11.105 65.515 11.275 ;
      LAYER via2 ;
        RECT 65.33 0.92 65.53 1.12 ;
    END
  END out[4]
  PIN out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 78.315 15.695 78.485 17.905 ;
        RECT 75.795 17.255 78.485 17.425 ;
        RECT 78.23 16.545 78.485 17.425 ;
        RECT 75.795 16.545 78.485 16.715 ;
        RECT 77.475 17.255 77.645 17.905 ;
        RECT 77.475 15.695 77.645 16.715 ;
        RECT 76.635 17.255 76.805 17.905 ;
        RECT 76.635 15.695 76.805 16.715 ;
        RECT 75.795 17.255 75.965 17.905 ;
        RECT 75.795 15.695 75.965 16.715 ;
      LAYER met1 ;
        RECT 76.31 16.5 76.63 16.76 ;
      LAYER met4 ;
        RECT 74.235 3.295 74.565 3.625 ;
        RECT 74.25 0 74.55 3.625 ;
      LAYER met3 ;
        RECT 76.305 3.295 76.635 3.625 ;
        RECT 74.21 3.31 76.635 3.61 ;
        RECT 74.21 3.3 74.59 3.62 ;
      LAYER met2 ;
        RECT 76.33 3.275 76.61 3.645 ;
        RECT 76.34 16.47 76.6 16.79 ;
        RECT 76.4 3.275 76.54 16.79 ;
      LAYER via3 ;
        RECT 74.3 3.36 74.5 3.56 ;
      LAYER via ;
        RECT 76.395 16.555 76.545 16.705 ;
      LAYER mcon ;
        RECT 76.385 16.545 76.555 16.715 ;
      LAYER via2 ;
        RECT 76.37 3.36 76.57 3.56 ;
    END
  END out[5]
  PIN out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 87.055 10.255 87.225 12.465 ;
        RECT 84.535 11.815 87.225 11.985 ;
        RECT 86.97 11.105 87.225 11.985 ;
        RECT 84.535 11.105 87.225 11.275 ;
        RECT 86.215 11.815 86.385 12.465 ;
        RECT 86.215 10.255 86.385 11.275 ;
        RECT 85.375 11.815 85.545 12.465 ;
        RECT 85.375 10.255 85.545 11.275 ;
        RECT 84.535 11.815 84.705 12.465 ;
        RECT 84.535 10.255 84.705 11.275 ;
      LAYER met1 ;
        RECT 87.35 10.38 87.67 10.64 ;
        RECT 86.905 11.12 87.58 11.26 ;
        RECT 87.44 10.38 87.58 11.26 ;
        RECT 86.905 11.075 87.195 11.305 ;
      LAYER met4 ;
        RECT 87.345 10.005 87.675 10.335 ;
        RECT 87.36 0 87.66 10.335 ;
      LAYER met3 ;
        RECT 87.32 10.01 87.7 10.33 ;
        RECT 87.345 10.005 87.675 10.335 ;
        RECT 86.9 10.02 87.7 10.32 ;
      LAYER met2 ;
        RECT 87.37 9.985 87.65 10.355 ;
        RECT 87.38 9.985 87.64 10.67 ;
      LAYER via3 ;
        RECT 87.41 10.07 87.61 10.27 ;
      LAYER via ;
        RECT 87.435 10.435 87.585 10.585 ;
      LAYER mcon ;
        RECT 86.965 11.105 87.135 11.275 ;
      LAYER via2 ;
        RECT 87.41 10.07 87.61 10.27 ;
    END
  END out[6]
  PIN out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 107.755 15.695 107.925 17.905 ;
        RECT 105.235 17.255 107.925 17.425 ;
        RECT 107.67 16.545 107.925 17.425 ;
        RECT 105.235 16.545 107.925 16.715 ;
        RECT 106.915 17.255 107.085 17.905 ;
        RECT 106.915 15.695 107.085 16.715 ;
        RECT 106.075 17.255 106.245 17.905 ;
        RECT 106.075 15.695 106.245 16.715 ;
        RECT 105.235 17.255 105.405 17.905 ;
        RECT 105.235 15.695 105.405 16.715 ;
      LAYER met1 ;
        RECT 105.305 16.515 105.595 16.745 ;
        RECT 105.38 16.22 105.52 16.745 ;
        RECT 101.15 16.22 105.52 16.36 ;
        RECT 101.15 16.16 101.47 16.42 ;
      LAYER met4 ;
        RECT 99.765 2.685 100.095 3.015 ;
        RECT 99.78 0 100.08 3.015 ;
      LAYER met3 ;
        RECT 101.145 2.685 101.475 3.015 ;
        RECT 99.74 2.7 101.475 3 ;
        RECT 99.74 2.69 100.12 3.01 ;
      LAYER met2 ;
        RECT 101.17 2.665 101.45 3.035 ;
        RECT 101.18 16.13 101.44 16.45 ;
        RECT 101.24 2.665 101.38 16.45 ;
      LAYER via3 ;
        RECT 99.83 2.75 100.03 2.95 ;
      LAYER via ;
        RECT 101.235 16.215 101.385 16.365 ;
      LAYER mcon ;
        RECT 105.365 16.545 105.535 16.715 ;
      LAYER via2 ;
        RECT 101.21 2.75 101.41 2.95 ;
    END
  END out[7]
  PIN out[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 112.855 19.605 113.025 20.625 ;
        RECT 110.335 18.895 113.025 19.065 ;
        RECT 112.855 18.415 113.025 19.065 ;
        RECT 110.335 19.605 113.025 19.775 ;
        RECT 112.015 19.605 112.185 20.625 ;
        RECT 112.015 18.415 112.185 19.065 ;
        RECT 111.175 19.605 111.345 20.625 ;
        RECT 111.175 18.415 111.345 19.065 ;
        RECT 110.335 18.895 110.595 19.095 ;
        RECT 110.335 18.895 110.59 19.775 ;
        RECT 110.335 18.415 110.505 20.625 ;
      LAYER met1 ;
        RECT 110.365 18.895 110.655 19.125 ;
        RECT 106.67 18.94 110.655 19.08 ;
        RECT 106.67 18.88 106.99 19.14 ;
      LAYER met4 ;
        RECT 112.875 8.785 113.205 9.115 ;
        RECT 112.89 0 113.19 9.115 ;
      LAYER met3 ;
        RECT 112.85 8.79 113.23 9.11 ;
        RECT 107.125 8.8 113.23 9.1 ;
        RECT 107.125 8.785 107.455 9.115 ;
      LAYER met2 ;
        RECT 107.15 8.765 107.43 9.135 ;
        RECT 106.76 9.76 107.36 9.9 ;
        RECT 107.22 8.765 107.36 9.9 ;
        RECT 106.7 18.85 106.96 19.17 ;
        RECT 106.76 9.76 106.9 19.17 ;
      LAYER via3 ;
        RECT 112.94 8.85 113.14 9.05 ;
      LAYER via ;
        RECT 106.755 18.935 106.905 19.085 ;
      LAYER mcon ;
        RECT 110.425 18.925 110.595 19.095 ;
      LAYER via2 ;
        RECT 107.19 8.85 107.39 9.05 ;
    END
  END out[8]
  PIN out[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 121.595 17.255 121.765 17.905 ;
        RECT 119.075 16.545 121.765 16.715 ;
        RECT 121.595 15.695 121.765 16.715 ;
        RECT 119.075 17.255 121.765 17.425 ;
        RECT 120.755 17.255 120.925 17.905 ;
        RECT 120.755 15.695 120.925 16.715 ;
        RECT 119.915 17.255 120.085 17.905 ;
        RECT 119.915 15.695 120.085 16.715 ;
        RECT 119.075 16.545 119.33 17.425 ;
        RECT 119.075 15.695 119.245 17.905 ;
      LAYER met1 ;
        RECT 120.47 16.5 120.79 16.76 ;
      LAYER met4 ;
        RECT 125.985 14.275 126.315 14.605 ;
        RECT 126 0 126.3 14.605 ;
      LAYER met3 ;
        RECT 125.96 14.28 126.34 14.6 ;
        RECT 120.465 14.29 126.34 14.59 ;
        RECT 120.465 14.275 120.795 14.605 ;
      LAYER met2 ;
        RECT 120.49 14.255 120.77 14.625 ;
        RECT 120.5 16.47 120.76 16.79 ;
        RECT 120.56 14.255 120.7 16.79 ;
      LAYER via3 ;
        RECT 126.05 14.34 126.25 14.54 ;
      LAYER via ;
        RECT 120.555 16.555 120.705 16.705 ;
      LAYER mcon ;
        RECT 120.545 16.545 120.715 16.715 ;
      LAYER via2 ;
        RECT 120.53 14.34 120.73 14.54 ;
    END
  END out[9]
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met5 ;
        RECT 0 24.3 200 26.3 ;
        RECT 0 44.7 200 46.7 ;
      LAYER li1 ;
        RECT 56.985 30.065 58.675 32.935 ;
        RECT 55.165 30.585 58.675 31.845 ;
        RECT 55.185 30.585 55.355 32.855 ;
        RECT 49.645 30.585 54.99 31.845 ;
        RECT 52.395 30.065 54.99 31.845 ;
        RECT 54.13 30.065 54.445 32.345 ;
        RECT 52.25 30.585 52.42 32.645 ;
        RECT 50.08 30.585 50.345 32.305 ;
        RECT 49.155 31.675 49.485 32.345 ;
        RECT 48.7 30.915 49.03 31.845 ;
        RECT 48.035 31.675 48.555 33.475 ;
        RECT 47.755 31.255 48.11 32.935 ;
        RECT 47.345 31.675 48.555 32.935 ;
        RECT 45.965 31.675 47.175 33.455 ;
        RECT 44.585 31.675 47.175 32.935 ;
        RECT 44.585 30.585 45.795 32.935 ;
        RECT 45.275 30.045 45.795 32.935 ;
        RECT 44.125 30.51 44.415 33.01 ;
        RECT 43.435 30.045 43.955 33.475 ;
        RECT 42.745 30.585 43.955 32.935 ;
        RECT 41.825 30.065 42.575 33.455 ;
        RECT 40.905 30.585 42.575 32.935 ;
        RECT 38.135 30.065 40.73 33.455 ;
        RECT 35.385 30.585 40.73 32.935 ;
        RECT 32.615 30.065 35.21 33.455 ;
        RECT 29.865 30.585 35.21 32.935 ;
        RECT 29.405 30.51 29.695 33.01 ;
        RECT 28.715 30.045 29.235 33.475 ;
        RECT 28.025 30.585 29.235 32.935 ;
        RECT 27.105 30.065 27.855 33.455 ;
        RECT 26.185 30.585 27.855 32.935 ;
        RECT 23.415 30.065 26.01 33.455 ;
        RECT 20.665 30.585 26.01 32.935 ;
        RECT 17.895 30.065 20.49 33.455 ;
        RECT 15.145 30.585 20.49 32.935 ;
        RECT 14.685 30.51 14.975 33.01 ;
        RECT 13.995 30.045 14.515 33.475 ;
        RECT 13.305 30.585 14.515 32.935 ;
        RECT 11.925 30.065 13.135 33.455 ;
        RECT 10.545 30.585 13.135 32.935 ;
        RECT 10 37.115 189.86 37.285 ;
        RECT 189.025 35.95 189.315 38.45 ;
        RECT 187.645 35.505 188.855 38.895 ;
        RECT 186.265 36.025 188.855 38.375 ;
        RECT 184.405 35.505 186.095 38.895 ;
        RECT 182.585 36.025 186.095 38.375 ;
        RECT 179.815 35.505 182.41 38.895 ;
        RECT 177.065 36.025 182.41 38.375 ;
        RECT 176.605 35.95 176.895 38.45 ;
        RECT 175.915 35.485 176.435 38.915 ;
        RECT 175.225 36.025 176.435 38.375 ;
        RECT 174.305 35.505 175.055 38.895 ;
        RECT 173.385 36.025 175.055 38.375 ;
        RECT 170.615 35.505 173.21 38.895 ;
        RECT 167.865 36.025 173.21 38.375 ;
        RECT 165.095 35.505 167.69 38.895 ;
        RECT 162.345 36.025 167.69 38.375 ;
        RECT 161.885 35.95 162.175 38.45 ;
        RECT 161.195 35.485 161.715 38.915 ;
        RECT 160.505 36.025 161.715 38.375 ;
        RECT 159.585 35.505 160.335 38.895 ;
        RECT 158.665 36.025 160.335 38.375 ;
        RECT 155.895 35.505 158.49 38.895 ;
        RECT 153.145 36.025 158.49 38.375 ;
        RECT 150.375 35.505 152.97 38.895 ;
        RECT 147.625 36.025 152.97 38.375 ;
        RECT 147.165 35.95 147.455 38.45 ;
        RECT 146.475 35.485 146.995 38.915 ;
        RECT 145.785 36.025 146.995 38.375 ;
        RECT 144.865 35.505 145.615 38.895 ;
        RECT 143.945 36.025 145.615 38.375 ;
        RECT 141.175 35.505 143.77 38.895 ;
        RECT 138.425 36.025 143.77 38.375 ;
        RECT 135.655 35.505 138.25 38.895 ;
        RECT 132.905 36.025 138.25 38.375 ;
        RECT 132.445 35.95 132.735 38.45 ;
        RECT 131.755 35.485 132.275 38.915 ;
        RECT 131.065 36.025 132.275 38.375 ;
        RECT 130.145 35.505 130.895 38.895 ;
        RECT 129.225 36.025 130.895 38.375 ;
        RECT 126.455 35.505 129.05 38.895 ;
        RECT 123.705 36.025 129.05 38.375 ;
        RECT 120.935 35.505 123.53 38.895 ;
        RECT 118.185 36.025 123.53 38.375 ;
        RECT 117.725 35.95 118.015 38.45 ;
        RECT 117.035 35.485 117.555 38.915 ;
        RECT 116.345 36.025 117.555 38.375 ;
        RECT 115.425 35.505 116.175 38.895 ;
        RECT 114.505 36.025 116.175 38.375 ;
        RECT 111.735 35.505 114.33 38.895 ;
        RECT 108.985 36.025 114.33 38.375 ;
        RECT 106.215 35.505 108.81 38.895 ;
        RECT 103.465 36.025 108.81 38.375 ;
        RECT 103.005 35.95 103.295 38.45 ;
        RECT 102.315 35.485 102.835 38.915 ;
        RECT 101.625 36.025 102.835 38.375 ;
        RECT 100.705 35.505 101.455 38.895 ;
        RECT 99.785 36.025 101.455 38.375 ;
        RECT 97.015 35.505 99.61 38.895 ;
        RECT 94.265 36.025 99.61 38.375 ;
        RECT 91.495 35.505 94.09 38.895 ;
        RECT 88.745 36.025 94.09 38.375 ;
        RECT 88.285 35.95 88.575 38.45 ;
        RECT 87.595 35.485 88.115 38.915 ;
        RECT 86.905 36.025 88.115 38.375 ;
        RECT 85.985 35.505 86.735 38.895 ;
        RECT 85.065 36.025 86.735 38.375 ;
        RECT 82.295 35.505 84.89 38.895 ;
        RECT 79.545 36.025 84.89 38.375 ;
        RECT 76.775 35.505 79.37 38.895 ;
        RECT 74.025 36.025 79.37 38.375 ;
        RECT 73.565 35.95 73.855 38.45 ;
        RECT 72.875 35.485 73.395 38.915 ;
        RECT 72.185 36.025 73.395 38.375 ;
        RECT 71.265 35.505 72.015 38.895 ;
        RECT 70.345 36.025 72.015 38.375 ;
        RECT 67.575 35.505 70.17 38.895 ;
        RECT 64.825 36.025 70.17 38.375 ;
        RECT 62.055 35.505 64.65 38.895 ;
        RECT 59.305 36.025 64.65 38.375 ;
        RECT 58.845 35.95 59.135 38.45 ;
        RECT 58.155 35.485 58.675 38.915 ;
        RECT 57.465 36.025 58.675 38.375 ;
        RECT 56.545 35.505 57.295 38.895 ;
        RECT 55.625 36.025 57.295 38.375 ;
        RECT 52.855 37.115 55.45 38.895 ;
        RECT 54.725 36.105 54.895 38.895 ;
        RECT 53.67 36.615 53.985 38.895 ;
        RECT 50.105 37.115 55.45 38.375 ;
        RECT 51.79 36.315 51.96 38.375 ;
        RECT 47.335 37.115 49.93 38.895 ;
        RECT 49.62 36.655 49.885 38.895 ;
        RECT 48.695 36.615 49.025 38.895 ;
        RECT 44.585 36.025 48.095 38.375 ;
        RECT 46.405 35.505 48.095 38.375 ;
        RECT 44.125 35.95 44.415 38.45 ;
        RECT 43.435 35.485 43.955 38.915 ;
        RECT 42.745 36.025 43.955 38.375 ;
        RECT 41.825 35.505 42.575 38.895 ;
        RECT 40.905 36.025 42.575 38.375 ;
        RECT 38.135 35.505 40.73 38.895 ;
        RECT 35.385 36.025 40.73 38.375 ;
        RECT 32.615 35.505 35.21 38.895 ;
        RECT 29.865 36.025 35.21 38.375 ;
        RECT 29.405 35.95 29.695 38.45 ;
        RECT 28.715 35.485 29.235 38.915 ;
        RECT 28.025 36.025 29.235 38.375 ;
        RECT 27.105 35.505 27.855 38.895 ;
        RECT 26.185 36.025 27.855 38.375 ;
        RECT 23.415 35.505 26.01 38.895 ;
        RECT 20.665 36.025 26.01 38.375 ;
        RECT 17.895 35.505 20.49 38.895 ;
        RECT 15.145 36.025 20.49 38.375 ;
        RECT 14.685 35.95 14.975 38.45 ;
        RECT 13.995 35.485 14.515 38.915 ;
        RECT 13.305 36.025 14.515 38.375 ;
        RECT 11.925 35.505 13.135 38.895 ;
        RECT 10.545 36.025 13.135 38.375 ;
        RECT 10 42.555 189.86 42.725 ;
        RECT 189.025 41.39 189.315 43.89 ;
        RECT 187.645 40.945 188.855 44.335 ;
        RECT 186.265 41.465 188.855 43.815 ;
        RECT 184.405 40.945 186.095 44.335 ;
        RECT 182.585 41.465 186.095 43.815 ;
        RECT 179.815 40.945 182.41 44.335 ;
        RECT 177.065 41.465 182.41 43.815 ;
        RECT 176.605 41.39 176.895 43.89 ;
        RECT 175.915 40.925 176.435 44.355 ;
        RECT 175.225 41.465 176.435 43.815 ;
        RECT 174.305 40.945 175.055 44.335 ;
        RECT 173.385 41.465 175.055 43.815 ;
        RECT 170.615 40.945 173.21 44.335 ;
        RECT 167.865 41.465 173.21 43.815 ;
        RECT 165.095 40.945 167.69 44.335 ;
        RECT 162.345 41.465 167.69 43.815 ;
        RECT 161.885 41.39 162.175 43.89 ;
        RECT 161.195 40.925 161.715 44.355 ;
        RECT 160.505 41.465 161.715 43.815 ;
        RECT 159.585 40.945 160.335 44.335 ;
        RECT 158.665 41.465 160.335 43.815 ;
        RECT 155.895 40.945 158.49 44.335 ;
        RECT 153.145 41.465 158.49 43.815 ;
        RECT 150.375 40.945 152.97 44.335 ;
        RECT 147.625 41.465 152.97 43.815 ;
        RECT 147.165 41.39 147.455 43.89 ;
        RECT 146.475 40.925 146.995 44.355 ;
        RECT 145.785 41.465 146.995 43.815 ;
        RECT 144.865 40.945 145.615 44.335 ;
        RECT 143.945 41.465 145.615 43.815 ;
        RECT 141.175 40.945 143.77 44.335 ;
        RECT 138.425 41.465 143.77 43.815 ;
        RECT 135.655 40.945 138.25 44.335 ;
        RECT 132.905 41.465 138.25 43.815 ;
        RECT 132.445 41.39 132.735 43.89 ;
        RECT 131.755 40.925 132.275 44.355 ;
        RECT 131.065 41.465 132.275 43.815 ;
        RECT 130.145 40.945 130.895 44.335 ;
        RECT 129.225 41.465 130.895 43.815 ;
        RECT 126.455 40.945 129.05 44.335 ;
        RECT 123.705 41.465 129.05 43.815 ;
        RECT 120.935 40.945 123.53 44.335 ;
        RECT 118.185 41.465 123.53 43.815 ;
        RECT 117.725 41.39 118.015 43.89 ;
        RECT 117.035 40.925 117.555 44.355 ;
        RECT 116.345 41.465 117.555 43.815 ;
        RECT 115.425 40.945 116.175 44.335 ;
        RECT 114.505 41.465 116.175 43.815 ;
        RECT 111.735 40.945 114.33 44.335 ;
        RECT 108.985 41.465 114.33 43.815 ;
        RECT 106.215 40.945 108.81 44.335 ;
        RECT 103.465 41.465 108.81 43.815 ;
        RECT 103.005 41.39 103.295 43.89 ;
        RECT 102.315 40.925 102.835 44.355 ;
        RECT 101.625 41.465 102.835 43.815 ;
        RECT 100.705 40.945 101.455 44.335 ;
        RECT 99.785 41.465 101.455 43.815 ;
        RECT 97.015 40.945 99.61 44.335 ;
        RECT 94.265 41.465 99.61 43.815 ;
        RECT 91.495 40.945 94.09 44.335 ;
        RECT 88.745 41.465 94.09 43.815 ;
        RECT 88.285 41.39 88.575 43.89 ;
        RECT 87.595 40.925 88.115 44.355 ;
        RECT 86.905 41.465 88.115 43.815 ;
        RECT 85.985 40.945 86.735 44.335 ;
        RECT 85.065 41.465 86.735 43.815 ;
        RECT 82.295 40.945 84.89 44.335 ;
        RECT 79.545 41.465 84.89 43.815 ;
        RECT 76.775 40.945 79.37 44.335 ;
        RECT 74.025 41.465 79.37 43.815 ;
        RECT 73.565 41.39 73.855 43.89 ;
        RECT 72.875 40.925 73.395 44.355 ;
        RECT 72.185 41.465 73.395 43.815 ;
        RECT 71.265 40.945 72.015 44.335 ;
        RECT 70.345 41.465 72.015 43.815 ;
        RECT 67.575 40.945 70.17 44.335 ;
        RECT 64.825 41.465 70.17 43.815 ;
        RECT 62.055 40.945 64.65 44.335 ;
        RECT 59.305 41.465 64.65 43.815 ;
        RECT 58.845 41.39 59.135 43.89 ;
        RECT 58.155 40.925 58.675 44.355 ;
        RECT 57.465 41.465 58.675 43.815 ;
        RECT 56.545 40.945 57.295 44.335 ;
        RECT 55.625 41.465 57.295 43.815 ;
        RECT 52.855 40.945 55.45 44.335 ;
        RECT 50.105 41.465 55.45 43.815 ;
        RECT 47.335 40.945 49.93 44.335 ;
        RECT 44.585 41.465 49.93 43.815 ;
        RECT 44.125 41.39 44.415 43.89 ;
        RECT 43.435 40.925 43.955 44.355 ;
        RECT 42.745 41.465 43.955 43.815 ;
        RECT 41.825 40.945 42.575 44.335 ;
        RECT 40.905 41.465 42.575 43.815 ;
        RECT 38.135 40.945 40.73 44.335 ;
        RECT 35.385 41.465 40.73 43.815 ;
        RECT 32.615 40.945 35.21 44.335 ;
        RECT 29.865 41.465 35.21 43.815 ;
        RECT 29.405 41.39 29.695 43.89 ;
        RECT 28.715 40.925 29.235 44.355 ;
        RECT 28.025 41.465 29.235 43.815 ;
        RECT 27.105 40.945 27.855 44.335 ;
        RECT 26.185 41.465 27.855 43.815 ;
        RECT 23.415 40.945 26.01 44.335 ;
        RECT 20.665 41.465 26.01 43.815 ;
        RECT 17.895 40.945 20.49 44.335 ;
        RECT 15.145 41.465 20.49 43.815 ;
        RECT 14.685 41.39 14.975 43.89 ;
        RECT 13.995 40.925 14.515 44.355 ;
        RECT 13.305 41.465 14.515 43.815 ;
        RECT 11.925 40.945 13.135 44.335 ;
        RECT 10.545 41.465 13.135 43.815 ;
        RECT 10 47.995 189.86 48.165 ;
        RECT 189.025 46.83 189.315 49.33 ;
        RECT 187.645 46.385 188.855 49.775 ;
        RECT 186.265 46.905 188.855 49.255 ;
        RECT 184.405 46.385 186.095 49.775 ;
        RECT 182.585 46.905 186.095 49.255 ;
        RECT 179.815 46.385 182.41 49.775 ;
        RECT 177.065 46.905 182.41 49.255 ;
        RECT 176.605 46.83 176.895 49.33 ;
        RECT 175.915 46.365 176.435 49.795 ;
        RECT 175.225 46.905 176.435 49.255 ;
        RECT 174.305 46.385 175.055 49.775 ;
        RECT 173.385 46.905 175.055 49.255 ;
        RECT 170.615 46.385 173.21 49.775 ;
        RECT 167.865 46.905 173.21 49.255 ;
        RECT 165.095 46.385 167.69 49.775 ;
        RECT 162.345 46.905 167.69 49.255 ;
        RECT 161.885 46.83 162.175 49.33 ;
        RECT 161.195 46.365 161.715 49.795 ;
        RECT 160.505 46.905 161.715 49.255 ;
        RECT 159.585 46.385 160.335 49.775 ;
        RECT 158.665 46.905 160.335 49.255 ;
        RECT 155.895 46.385 158.49 49.775 ;
        RECT 153.145 46.905 158.49 49.255 ;
        RECT 150.375 46.385 152.97 49.775 ;
        RECT 147.625 46.905 152.97 49.255 ;
        RECT 147.165 46.83 147.455 49.33 ;
        RECT 146.475 46.365 146.995 49.795 ;
        RECT 145.785 46.905 146.995 49.255 ;
        RECT 144.865 46.385 145.615 49.775 ;
        RECT 143.945 46.905 145.615 49.255 ;
        RECT 141.175 46.385 143.77 49.775 ;
        RECT 138.425 46.905 143.77 49.255 ;
        RECT 135.655 46.385 138.25 49.775 ;
        RECT 132.905 46.905 138.25 49.255 ;
        RECT 132.445 46.83 132.735 49.33 ;
        RECT 131.755 46.365 132.275 49.795 ;
        RECT 131.065 46.905 132.275 49.255 ;
        RECT 130.145 46.385 130.895 49.775 ;
        RECT 129.225 46.905 130.895 49.255 ;
        RECT 126.455 46.385 129.05 49.775 ;
        RECT 123.705 46.905 129.05 49.255 ;
        RECT 120.935 46.385 123.53 49.775 ;
        RECT 118.185 46.905 123.53 49.255 ;
        RECT 117.725 46.83 118.015 49.33 ;
        RECT 117.035 46.365 117.555 49.795 ;
        RECT 116.345 46.905 117.555 49.255 ;
        RECT 115.425 46.385 116.175 49.775 ;
        RECT 114.505 46.905 116.175 49.255 ;
        RECT 111.735 46.385 114.33 49.775 ;
        RECT 108.985 46.905 114.33 49.255 ;
        RECT 106.215 46.385 108.81 49.775 ;
        RECT 103.465 46.905 108.81 49.255 ;
        RECT 103.005 46.83 103.295 49.33 ;
        RECT 102.315 46.365 102.835 49.795 ;
        RECT 101.625 46.905 102.835 49.255 ;
        RECT 100.705 46.385 101.455 49.775 ;
        RECT 99.785 46.905 101.455 49.255 ;
        RECT 97.015 46.385 99.61 49.775 ;
        RECT 94.265 46.905 99.61 49.255 ;
        RECT 91.495 46.385 94.09 49.775 ;
        RECT 88.745 46.905 94.09 49.255 ;
        RECT 88.285 46.83 88.575 49.33 ;
        RECT 87.595 46.365 88.115 49.795 ;
        RECT 86.905 46.905 88.115 49.255 ;
        RECT 85.985 46.385 86.735 49.775 ;
        RECT 85.065 46.905 86.735 49.255 ;
        RECT 82.295 46.385 84.89 49.775 ;
        RECT 79.545 46.905 84.89 49.255 ;
        RECT 76.775 46.385 79.37 49.775 ;
        RECT 74.025 46.905 79.37 49.255 ;
        RECT 73.565 46.83 73.855 49.33 ;
        RECT 72.875 46.365 73.395 49.795 ;
        RECT 72.185 46.905 73.395 49.255 ;
        RECT 71.265 46.385 72.015 49.775 ;
        RECT 70.345 46.905 72.015 49.255 ;
        RECT 67.575 46.385 70.17 49.775 ;
        RECT 64.825 46.905 70.17 49.255 ;
        RECT 62.055 46.385 64.65 49.775 ;
        RECT 59.305 46.905 64.65 49.255 ;
        RECT 58.845 46.83 59.135 49.33 ;
        RECT 58.155 46.365 58.675 49.795 ;
        RECT 57.465 46.905 58.675 49.255 ;
        RECT 56.545 46.385 57.295 49.775 ;
        RECT 55.625 46.905 57.295 49.255 ;
        RECT 52.855 46.385 55.45 49.775 ;
        RECT 50.105 46.905 55.45 49.255 ;
        RECT 47.335 46.385 49.93 49.775 ;
        RECT 44.585 46.905 49.93 49.255 ;
        RECT 44.125 46.83 44.415 49.33 ;
        RECT 43.435 46.365 43.955 49.795 ;
        RECT 42.745 46.905 43.955 49.255 ;
        RECT 41.825 46.385 42.575 49.775 ;
        RECT 40.905 46.905 42.575 49.255 ;
        RECT 38.135 46.385 40.73 49.775 ;
        RECT 35.385 46.905 40.73 49.255 ;
        RECT 32.615 46.385 35.21 49.775 ;
        RECT 29.865 46.905 35.21 49.255 ;
        RECT 29.405 46.83 29.695 49.33 ;
        RECT 28.715 46.365 29.235 49.795 ;
        RECT 28.025 46.905 29.235 49.255 ;
        RECT 27.105 46.385 27.855 49.775 ;
        RECT 26.185 46.905 27.855 49.255 ;
        RECT 23.415 46.385 26.01 49.775 ;
        RECT 20.665 46.905 26.01 49.255 ;
        RECT 17.895 46.385 20.49 49.775 ;
        RECT 15.145 46.905 20.49 49.255 ;
        RECT 14.685 46.83 14.975 49.33 ;
        RECT 13.995 46.365 14.515 49.795 ;
        RECT 13.305 46.905 14.515 49.255 ;
        RECT 11.925 46.385 13.135 49.775 ;
        RECT 10.545 46.905 13.135 49.255 ;
        RECT 10 53.435 189.86 53.605 ;
        RECT 189.025 52.27 189.315 54.77 ;
        RECT 187.645 51.825 188.855 55.215 ;
        RECT 186.265 52.345 188.855 54.695 ;
        RECT 184.405 51.825 186.095 55.215 ;
        RECT 182.585 52.345 186.095 54.695 ;
        RECT 179.815 51.825 182.41 55.215 ;
        RECT 177.065 52.345 182.41 54.695 ;
        RECT 176.605 52.27 176.895 54.77 ;
        RECT 175.915 51.805 176.435 55.235 ;
        RECT 175.225 52.345 176.435 54.695 ;
        RECT 174.305 51.825 175.055 55.215 ;
        RECT 173.385 52.345 175.055 54.695 ;
        RECT 170.615 51.825 173.21 55.215 ;
        RECT 167.865 52.345 173.21 54.695 ;
        RECT 165.095 51.825 167.69 55.215 ;
        RECT 162.345 52.345 167.69 54.695 ;
        RECT 161.885 52.27 162.175 54.77 ;
        RECT 161.195 51.805 161.715 55.235 ;
        RECT 160.505 52.345 161.715 54.695 ;
        RECT 159.585 51.825 160.335 55.215 ;
        RECT 158.665 52.345 160.335 54.695 ;
        RECT 155.895 51.825 158.49 55.215 ;
        RECT 153.145 52.345 158.49 54.695 ;
        RECT 150.375 51.825 152.97 55.215 ;
        RECT 147.625 52.345 152.97 54.695 ;
        RECT 147.165 52.27 147.455 54.77 ;
        RECT 146.475 51.805 146.995 55.235 ;
        RECT 145.785 52.345 146.995 54.695 ;
        RECT 144.865 51.825 145.615 55.215 ;
        RECT 143.945 52.345 145.615 54.695 ;
        RECT 141.175 51.825 143.77 55.215 ;
        RECT 138.425 52.345 143.77 54.695 ;
        RECT 135.655 51.825 138.25 55.215 ;
        RECT 132.905 52.345 138.25 54.695 ;
        RECT 132.445 52.27 132.735 54.77 ;
        RECT 131.755 51.805 132.275 55.235 ;
        RECT 131.065 52.345 132.275 54.695 ;
        RECT 130.145 51.825 130.895 55.215 ;
        RECT 129.225 52.345 130.895 54.695 ;
        RECT 126.455 51.825 129.05 55.215 ;
        RECT 123.705 52.345 129.05 54.695 ;
        RECT 120.935 51.825 123.53 55.215 ;
        RECT 118.185 52.345 123.53 54.695 ;
        RECT 117.725 52.27 118.015 54.77 ;
        RECT 117.035 51.805 117.555 55.235 ;
        RECT 116.345 52.345 117.555 54.695 ;
        RECT 115.425 51.825 116.175 55.215 ;
        RECT 114.505 52.345 116.175 54.695 ;
        RECT 111.735 51.825 114.33 55.215 ;
        RECT 108.985 52.345 114.33 54.695 ;
        RECT 106.215 51.825 108.81 55.215 ;
        RECT 103.465 52.345 108.81 54.695 ;
        RECT 103.005 52.27 103.295 54.77 ;
        RECT 102.315 51.805 102.835 55.235 ;
        RECT 101.625 52.345 102.835 54.695 ;
        RECT 100.705 51.825 101.455 55.215 ;
        RECT 99.785 52.345 101.455 54.695 ;
        RECT 97.015 51.825 99.61 55.215 ;
        RECT 94.265 52.345 99.61 54.695 ;
        RECT 91.495 51.825 94.09 55.215 ;
        RECT 88.745 52.345 94.09 54.695 ;
        RECT 88.285 52.27 88.575 54.77 ;
        RECT 87.595 51.805 88.115 55.235 ;
        RECT 86.905 52.345 88.115 54.695 ;
        RECT 85.985 51.825 86.735 55.215 ;
        RECT 85.065 52.345 86.735 54.695 ;
        RECT 82.295 51.825 84.89 55.215 ;
        RECT 79.545 52.345 84.89 54.695 ;
        RECT 76.775 51.825 79.37 55.215 ;
        RECT 74.025 52.345 79.37 54.695 ;
        RECT 73.565 52.27 73.855 54.77 ;
        RECT 72.875 51.805 73.395 55.235 ;
        RECT 72.185 52.345 73.395 54.695 ;
        RECT 71.265 51.825 72.015 55.215 ;
        RECT 70.345 52.345 72.015 54.695 ;
        RECT 67.575 51.825 70.17 55.215 ;
        RECT 64.825 52.345 70.17 54.695 ;
        RECT 62.055 51.825 64.65 55.215 ;
        RECT 59.305 52.345 64.65 54.695 ;
        RECT 58.845 52.27 59.135 54.77 ;
        RECT 58.155 51.805 58.675 55.235 ;
        RECT 57.465 52.345 58.675 54.695 ;
        RECT 56.545 51.825 57.295 55.215 ;
        RECT 55.625 52.345 57.295 54.695 ;
        RECT 52.855 51.825 55.45 55.215 ;
        RECT 50.105 52.345 55.45 54.695 ;
        RECT 47.335 51.825 49.93 55.215 ;
        RECT 44.585 52.345 49.93 54.695 ;
        RECT 44.125 52.27 44.415 54.77 ;
        RECT 43.435 51.805 43.955 55.235 ;
        RECT 42.745 52.345 43.955 54.695 ;
        RECT 41.825 51.825 42.575 55.215 ;
        RECT 40.905 52.345 42.575 54.695 ;
        RECT 38.135 51.825 40.73 55.215 ;
        RECT 35.385 52.345 40.73 54.695 ;
        RECT 32.615 51.825 35.21 55.215 ;
        RECT 29.865 52.345 35.21 54.695 ;
        RECT 29.405 52.27 29.695 54.77 ;
        RECT 28.715 51.805 29.235 55.235 ;
        RECT 28.025 52.345 29.235 54.695 ;
        RECT 27.105 51.825 27.855 55.215 ;
        RECT 26.185 52.345 27.855 54.695 ;
        RECT 23.415 51.825 26.01 55.215 ;
        RECT 20.665 52.345 26.01 54.695 ;
        RECT 17.895 51.825 20.49 55.215 ;
        RECT 15.145 52.345 20.49 54.695 ;
        RECT 14.685 52.27 14.975 54.77 ;
        RECT 13.995 51.805 14.515 55.235 ;
        RECT 13.305 52.345 14.515 54.695 ;
        RECT 11.925 51.825 13.135 55.215 ;
        RECT 10.545 52.345 13.135 54.695 ;
        RECT 10 58.875 189.86 59.045 ;
        RECT 189.025 57.71 189.315 59.045 ;
        RECT 186.265 57.785 188.855 59.045 ;
        RECT 187.645 57.265 188.855 59.045 ;
        RECT 182.585 57.785 186.095 59.045 ;
        RECT 184.405 57.265 186.095 59.045 ;
        RECT 177.065 57.785 182.41 59.045 ;
        RECT 179.815 57.265 182.41 59.045 ;
        RECT 176.605 57.71 176.895 59.045 ;
        RECT 175.225 57.785 176.435 59.045 ;
        RECT 175.915 57.245 176.435 59.045 ;
        RECT 173.385 57.785 175.055 59.045 ;
        RECT 174.305 57.265 175.055 59.045 ;
        RECT 167.865 57.785 173.21 59.045 ;
        RECT 170.615 57.265 173.21 59.045 ;
        RECT 162.345 57.785 167.69 59.045 ;
        RECT 165.095 57.265 167.69 59.045 ;
        RECT 161.885 57.71 162.175 59.045 ;
        RECT 160.505 57.785 161.715 59.045 ;
        RECT 161.195 57.245 161.715 59.045 ;
        RECT 158.665 57.785 160.335 59.045 ;
        RECT 159.585 57.265 160.335 59.045 ;
        RECT 153.145 57.785 158.49 59.045 ;
        RECT 155.895 57.265 158.49 59.045 ;
        RECT 147.625 57.785 152.97 59.045 ;
        RECT 150.375 57.265 152.97 59.045 ;
        RECT 147.165 57.71 147.455 59.045 ;
        RECT 145.785 57.785 146.995 59.045 ;
        RECT 146.475 57.245 146.995 59.045 ;
        RECT 143.945 57.785 145.615 59.045 ;
        RECT 144.865 57.265 145.615 59.045 ;
        RECT 138.425 57.785 143.77 59.045 ;
        RECT 141.175 57.265 143.77 59.045 ;
        RECT 132.905 57.785 138.25 59.045 ;
        RECT 135.655 57.265 138.25 59.045 ;
        RECT 132.445 57.71 132.735 59.045 ;
        RECT 131.065 57.785 132.275 59.045 ;
        RECT 131.755 57.245 132.275 59.045 ;
        RECT 129.225 57.785 130.895 59.045 ;
        RECT 130.145 57.265 130.895 59.045 ;
        RECT 123.705 57.785 129.05 59.045 ;
        RECT 126.455 57.265 129.05 59.045 ;
        RECT 118.185 57.785 123.53 59.045 ;
        RECT 120.935 57.265 123.53 59.045 ;
        RECT 117.725 57.71 118.015 59.045 ;
        RECT 116.345 57.785 117.555 59.045 ;
        RECT 117.035 57.245 117.555 59.045 ;
        RECT 114.505 57.785 116.175 59.045 ;
        RECT 115.425 57.265 116.175 59.045 ;
        RECT 108.985 57.785 114.33 59.045 ;
        RECT 111.735 57.265 114.33 59.045 ;
        RECT 103.465 57.785 108.81 59.045 ;
        RECT 106.215 57.265 108.81 59.045 ;
        RECT 103.005 57.71 103.295 59.045 ;
        RECT 101.625 57.785 102.835 59.045 ;
        RECT 102.315 57.245 102.835 59.045 ;
        RECT 99.785 57.785 101.455 59.045 ;
        RECT 100.705 57.265 101.455 59.045 ;
        RECT 94.265 57.785 99.61 59.045 ;
        RECT 97.015 57.265 99.61 59.045 ;
        RECT 88.745 57.785 94.09 59.045 ;
        RECT 91.495 57.265 94.09 59.045 ;
        RECT 88.285 57.71 88.575 59.045 ;
        RECT 86.905 57.785 88.115 59.045 ;
        RECT 87.595 57.245 88.115 59.045 ;
        RECT 85.065 57.785 86.735 59.045 ;
        RECT 85.985 57.265 86.735 59.045 ;
        RECT 79.545 57.785 84.89 59.045 ;
        RECT 82.295 57.265 84.89 59.045 ;
        RECT 74.025 57.785 79.37 59.045 ;
        RECT 76.775 57.265 79.37 59.045 ;
        RECT 73.565 57.71 73.855 59.045 ;
        RECT 72.185 57.785 73.395 59.045 ;
        RECT 72.875 57.245 73.395 59.045 ;
        RECT 70.345 57.785 72.015 59.045 ;
        RECT 71.265 57.265 72.015 59.045 ;
        RECT 64.825 57.785 70.17 59.045 ;
        RECT 67.575 57.265 70.17 59.045 ;
        RECT 59.305 57.785 64.65 59.045 ;
        RECT 62.055 57.265 64.65 59.045 ;
        RECT 58.845 57.71 59.135 59.045 ;
        RECT 57.465 57.785 58.675 59.045 ;
        RECT 58.155 57.245 58.675 59.045 ;
        RECT 55.625 57.785 57.295 59.045 ;
        RECT 56.545 57.265 57.295 59.045 ;
        RECT 50.105 57.785 55.45 59.045 ;
        RECT 52.855 57.265 55.45 59.045 ;
        RECT 44.585 57.785 49.93 59.045 ;
        RECT 47.335 57.265 49.93 59.045 ;
        RECT 44.125 57.71 44.415 59.045 ;
        RECT 42.745 57.785 43.955 59.045 ;
        RECT 43.435 57.245 43.955 59.045 ;
        RECT 40.905 57.785 42.575 59.045 ;
        RECT 41.825 57.265 42.575 59.045 ;
        RECT 35.385 57.785 40.73 59.045 ;
        RECT 38.135 57.265 40.73 59.045 ;
        RECT 29.865 57.785 35.21 59.045 ;
        RECT 32.615 57.265 35.21 59.045 ;
        RECT 29.405 57.71 29.695 59.045 ;
        RECT 28.025 57.785 29.235 59.045 ;
        RECT 28.715 57.245 29.235 59.045 ;
        RECT 26.185 57.785 27.855 59.045 ;
        RECT 27.105 57.265 27.855 59.045 ;
        RECT 20.665 57.785 26.01 59.045 ;
        RECT 23.415 57.265 26.01 59.045 ;
        RECT 15.145 57.785 20.49 59.045 ;
        RECT 17.895 57.265 20.49 59.045 ;
        RECT 14.685 57.71 14.975 59.045 ;
        RECT 13.305 57.785 14.515 59.045 ;
        RECT 13.995 57.245 14.515 59.045 ;
        RECT 10.545 57.785 13.135 59.045 ;
        RECT 11.925 57.265 13.135 59.045 ;
        RECT 10 9.915 189.86 10.085 ;
        RECT 189.025 9.915 189.315 11.25 ;
        RECT 187.645 9.915 188.855 11.695 ;
        RECT 186.265 9.915 188.855 11.175 ;
        RECT 184.405 9.915 186.095 11.695 ;
        RECT 182.585 9.915 186.095 11.175 ;
        RECT 179.815 9.915 182.41 11.695 ;
        RECT 177.065 9.915 182.41 11.175 ;
        RECT 176.605 9.915 176.895 11.25 ;
        RECT 175.915 9.915 176.435 11.715 ;
        RECT 175.225 9.915 176.435 11.175 ;
        RECT 173.845 9.915 175.055 11.695 ;
        RECT 172.465 9.915 175.055 11.175 ;
        RECT 170.605 9.915 172.295 11.695 ;
        RECT 168.785 9.915 172.295 11.175 ;
        RECT 167.895 9.915 168.225 11.235 ;
        RECT 167.055 9.915 167.385 10.885 ;
        RECT 166.215 9.915 166.545 10.885 ;
        RECT 165.375 9.915 165.705 10.885 ;
        RECT 164.615 9.915 164.785 10.885 ;
        RECT 163.775 9.915 163.945 10.885 ;
        RECT 161.885 9.915 162.175 11.25 ;
        RECT 161.195 9.915 161.715 11.715 ;
        RECT 160.505 9.915 161.715 11.175 ;
        RECT 159.125 9.915 160.335 11.695 ;
        RECT 157.745 9.915 160.335 11.175 ;
        RECT 155.885 9.915 157.575 11.695 ;
        RECT 154.065 9.915 157.575 11.175 ;
        RECT 153.175 9.915 153.505 11.235 ;
        RECT 152.335 9.915 152.665 10.885 ;
        RECT 151.495 9.915 151.825 10.885 ;
        RECT 150.655 9.915 150.985 10.885 ;
        RECT 149.895 9.915 150.065 10.885 ;
        RECT 149.055 9.915 149.225 10.885 ;
        RECT 147.165 9.915 147.455 11.25 ;
        RECT 146.475 9.915 146.995 11.715 ;
        RECT 145.785 9.915 146.995 11.175 ;
        RECT 144.865 9.915 145.615 11.695 ;
        RECT 143.945 9.915 145.615 11.175 ;
        RECT 143.055 9.915 143.385 11.235 ;
        RECT 142.215 9.915 142.545 10.885 ;
        RECT 141.375 9.915 141.705 10.885 ;
        RECT 140.535 9.915 140.865 10.885 ;
        RECT 139.775 9.915 139.945 10.885 ;
        RECT 138.935 9.915 139.105 10.885 ;
        RECT 135.655 9.915 138.25 11.695 ;
        RECT 132.905 9.915 138.25 11.175 ;
        RECT 132.445 9.915 132.735 11.25 ;
        RECT 131.755 9.915 132.275 11.715 ;
        RECT 131.065 9.915 132.275 11.175 ;
        RECT 130.145 9.915 130.895 11.695 ;
        RECT 129.225 9.915 130.895 11.175 ;
        RECT 126.455 9.915 129.05 11.695 ;
        RECT 123.705 9.915 129.05 11.175 ;
        RECT 122.855 9.915 123.025 10.885 ;
        RECT 122.015 9.915 122.185 10.885 ;
        RECT 121.095 9.915 121.425 10.885 ;
        RECT 120.255 9.915 120.585 10.885 ;
        RECT 119.415 9.915 119.745 10.885 ;
        RECT 118.575 9.915 118.905 11.235 ;
        RECT 117.725 9.915 118.015 11.25 ;
        RECT 117.035 9.915 117.555 11.715 ;
        RECT 116.345 9.915 117.555 11.175 ;
        RECT 115.425 9.915 116.175 11.695 ;
        RECT 114.505 9.915 116.175 11.175 ;
        RECT 111.735 9.915 114.33 11.695 ;
        RECT 108.985 9.915 114.33 11.175 ;
        RECT 106.215 9.915 108.81 11.695 ;
        RECT 103.465 9.915 108.81 11.175 ;
        RECT 103.005 9.915 103.295 11.25 ;
        RECT 102.115 9.915 102.445 11.235 ;
        RECT 101.275 9.915 101.605 10.885 ;
        RECT 100.435 9.915 100.765 10.885 ;
        RECT 99.595 9.915 99.925 10.885 ;
        RECT 98.835 9.915 99.005 10.885 ;
        RECT 97.995 9.915 98.165 10.885 ;
        RECT 96.135 9.915 96.465 11.235 ;
        RECT 95.295 9.915 95.625 10.885 ;
        RECT 94.455 9.915 94.785 10.885 ;
        RECT 93.615 9.915 93.945 10.885 ;
        RECT 92.855 9.915 93.025 10.885 ;
        RECT 92.015 9.915 92.185 10.885 ;
        RECT 90.125 9.915 91.335 11.695 ;
        RECT 88.745 9.915 91.335 11.175 ;
        RECT 88.285 9.915 88.575 11.25 ;
        RECT 87.395 9.915 87.725 11.235 ;
        RECT 86.555 9.915 86.885 10.885 ;
        RECT 85.715 9.915 86.045 10.885 ;
        RECT 84.875 9.915 85.205 10.885 ;
        RECT 84.115 9.915 84.285 10.885 ;
        RECT 83.275 9.915 83.445 10.885 ;
        RECT 82.075 9.915 82.595 11.715 ;
        RECT 81.385 9.915 82.595 11.175 ;
        RECT 80.465 9.915 81.215 11.695 ;
        RECT 79.545 9.915 81.215 11.175 ;
        RECT 78.655 9.915 78.985 11.235 ;
        RECT 77.815 9.915 78.145 10.885 ;
        RECT 76.975 9.915 77.305 10.885 ;
        RECT 76.135 9.915 76.465 10.885 ;
        RECT 75.375 9.915 75.545 10.885 ;
        RECT 74.535 9.915 74.705 10.885 ;
        RECT 73.565 9.915 73.855 11.25 ;
        RECT 70.795 9.915 73.39 11.695 ;
        RECT 68.045 9.915 73.39 11.175 ;
        RECT 67.155 9.915 67.485 11.235 ;
        RECT 66.315 9.915 66.645 10.885 ;
        RECT 65.475 9.915 65.805 10.885 ;
        RECT 64.635 9.915 64.965 10.885 ;
        RECT 63.875 9.915 64.045 10.885 ;
        RECT 63.035 9.915 63.205 10.885 ;
        RECT 61.835 9.915 62.355 11.715 ;
        RECT 61.145 9.915 62.355 11.175 ;
        RECT 60.225 9.915 60.975 11.695 ;
        RECT 59.305 9.915 60.975 11.175 ;
        RECT 58.845 9.915 59.135 11.25 ;
        RECT 56.075 9.915 58.67 11.695 ;
        RECT 53.325 9.915 58.67 11.175 ;
        RECT 52.435 9.915 52.765 11.235 ;
        RECT 51.595 9.915 51.925 10.885 ;
        RECT 50.755 9.915 51.085 10.885 ;
        RECT 49.915 9.915 50.245 10.885 ;
        RECT 49.155 9.915 49.325 10.885 ;
        RECT 48.315 9.915 48.485 10.885 ;
        RECT 47.115 9.915 47.635 11.715 ;
        RECT 46.425 9.915 47.635 11.175 ;
        RECT 45.505 9.915 46.255 11.695 ;
        RECT 44.585 9.915 46.255 11.175 ;
        RECT 44.125 9.915 44.415 11.25 ;
        RECT 43.435 9.915 43.955 11.715 ;
        RECT 42.745 9.915 43.955 11.175 ;
        RECT 41.825 9.915 42.575 11.695 ;
        RECT 40.905 9.915 42.575 11.175 ;
        RECT 38.135 9.915 40.73 11.695 ;
        RECT 35.385 9.915 40.73 11.175 ;
        RECT 34.495 9.915 34.825 11.235 ;
        RECT 33.655 9.915 33.985 10.885 ;
        RECT 32.815 9.915 33.145 10.885 ;
        RECT 31.975 9.915 32.305 10.885 ;
        RECT 31.215 9.915 31.385 10.885 ;
        RECT 30.375 9.915 30.545 10.885 ;
        RECT 29.405 9.915 29.695 11.25 ;
        RECT 28.715 9.915 29.235 11.715 ;
        RECT 28.025 9.915 29.235 11.175 ;
        RECT 27.105 9.915 27.855 11.695 ;
        RECT 26.185 9.915 27.855 11.175 ;
        RECT 23.415 9.915 26.01 11.695 ;
        RECT 20.665 9.915 26.01 11.175 ;
        RECT 17.895 9.915 20.49 11.695 ;
        RECT 15.145 9.915 20.49 11.175 ;
        RECT 14.685 9.915 14.975 11.25 ;
        RECT 13.995 9.915 14.515 11.715 ;
        RECT 13.305 9.915 14.515 11.175 ;
        RECT 11.925 9.915 13.135 11.695 ;
        RECT 10.545 9.915 13.135 11.175 ;
        RECT 10 15.355 189.86 15.525 ;
        RECT 189.025 14.19 189.315 16.69 ;
        RECT 187.645 13.745 188.855 17.135 ;
        RECT 186.265 14.265 188.855 16.615 ;
        RECT 184.405 13.745 186.095 17.135 ;
        RECT 182.585 14.265 186.095 16.615 ;
        RECT 177.065 14.265 182.41 15.525 ;
        RECT 179.815 13.745 182.41 15.525 ;
        RECT 181.695 13.745 182.025 16.675 ;
        RECT 180.855 13.745 181.185 16.325 ;
        RECT 180.015 13.745 180.345 16.325 ;
        RECT 179.175 14.265 179.505 16.325 ;
        RECT 178.415 14.265 178.585 16.325 ;
        RECT 177.575 14.265 177.745 16.325 ;
        RECT 176.605 14.19 176.895 16.69 ;
        RECT 175.225 14.265 176.435 15.525 ;
        RECT 175.915 13.725 176.435 15.525 ;
        RECT 175.705 14.265 175.875 16.535 ;
        RECT 171.545 14.265 175.055 15.525 ;
        RECT 173.365 13.745 175.055 15.525 ;
        RECT 174.65 13.745 174.965 16.025 ;
        RECT 172.77 14.265 172.94 16.325 ;
        RECT 170.6 15.355 170.865 15.985 ;
        RECT 169.675 15.355 170.005 16.025 ;
        RECT 169.23 14.935 169.585 15.525 ;
        RECT 168.555 15.355 169.075 17.155 ;
        RECT 168.31 14.595 168.64 16.615 ;
        RECT 167.865 15.355 169.075 16.615 ;
        RECT 162.345 14.265 167.69 15.525 ;
        RECT 165.095 13.745 167.69 15.525 ;
        RECT 166.975 13.745 167.305 16.675 ;
        RECT 166.135 13.745 166.465 16.325 ;
        RECT 165.295 13.745 165.625 16.325 ;
        RECT 164.455 14.265 164.785 16.325 ;
        RECT 163.695 14.265 163.865 16.325 ;
        RECT 162.855 14.265 163.025 16.325 ;
        RECT 161.885 14.19 162.175 16.69 ;
        RECT 160.505 14.265 161.715 15.525 ;
        RECT 161.195 13.725 161.715 15.525 ;
        RECT 158.665 14.265 160.335 15.525 ;
        RECT 159.585 13.745 160.335 15.525 ;
        RECT 160.065 13.745 160.235 16.535 ;
        RECT 159.01 14.265 159.325 16.025 ;
        RECT 153.145 14.265 158.49 15.525 ;
        RECT 155.895 13.745 158.49 15.525 ;
        RECT 157.13 13.745 157.3 16.325 ;
        RECT 154.96 14.265 155.225 15.985 ;
        RECT 154.035 14.265 154.365 16.025 ;
        RECT 152.915 15.355 153.435 17.155 ;
        RECT 147.625 14.265 152.97 15.525 ;
        RECT 152.225 15.355 153.435 16.615 ;
        RECT 150.375 13.745 152.97 15.525 ;
        RECT 151.305 13.745 152.055 17.135 ;
        RECT 150.385 13.745 152.055 16.615 ;
        RECT 149.005 14.265 150.215 17.135 ;
        RECT 147.625 14.265 150.215 16.615 ;
        RECT 147.165 14.19 147.455 16.69 ;
        RECT 144.865 14.265 146.075 15.525 ;
        RECT 145.555 13.725 146.075 15.525 ;
        RECT 145.3 14.265 145.63 16.285 ;
        RECT 144.355 15.355 144.71 15.945 ;
        RECT 144.015 14.555 144.185 15.525 ;
        RECT 143.175 14.555 143.345 15.525 ;
        RECT 142.255 14.555 142.585 15.525 ;
        RECT 141.875 15.355 142.395 17.155 ;
        RECT 141.185 15.355 142.395 16.615 ;
        RECT 141.415 14.555 141.745 16.615 ;
        RECT 139.805 15.355 141.015 17.135 ;
        RECT 140.575 14.555 140.905 17.135 ;
        RECT 139.735 14.205 140.065 16.615 ;
        RECT 138.425 15.355 141.015 16.615 ;
        RECT 137.535 14.205 137.865 15.525 ;
        RECT 137.48 15.355 137.81 16.285 ;
        RECT 136.695 14.555 137.025 15.525 ;
        RECT 136.535 15.355 136.89 15.945 ;
        RECT 135.855 14.555 136.185 15.525 ;
        RECT 135.015 14.555 135.345 15.525 ;
        RECT 133.825 15.355 134.575 17.135 ;
        RECT 134.255 14.555 134.425 17.135 ;
        RECT 132.905 15.355 134.575 16.615 ;
        RECT 133.415 14.555 133.585 16.615 ;
        RECT 132.445 14.19 132.735 16.69 ;
        RECT 131.755 13.725 132.275 17.155 ;
        RECT 131.065 14.265 132.275 16.615 ;
        RECT 130.145 13.745 130.895 17.135 ;
        RECT 129.225 13.745 130.895 16.615 ;
        RECT 127.385 14.265 130.895 15.525 ;
        RECT 129.205 13.745 130.895 15.525 ;
        RECT 128.28 14.265 128.61 16.285 ;
        RECT 127.335 15.355 127.69 15.945 ;
        RECT 121.865 14.265 127.21 15.525 ;
        RECT 124.615 13.745 127.21 15.525 ;
        RECT 124.625 13.745 125.375 17.135 ;
        RECT 123.705 14.265 125.375 16.615 ;
        RECT 122.855 14.265 123.025 16.325 ;
        RECT 122.015 14.265 122.185 16.325 ;
        RECT 121.095 15.355 121.425 16.325 ;
        RECT 120.92 14.595 121.25 15.525 ;
        RECT 120.255 15.355 120.585 16.325 ;
        RECT 119.975 14.935 120.33 15.525 ;
        RECT 119.415 15.355 119.745 16.325 ;
        RECT 118.575 15.355 118.905 16.675 ;
        RECT 117.725 14.19 118.015 16.69 ;
        RECT 116.345 14.265 117.555 17.135 ;
        RECT 116.805 13.745 117.555 17.135 ;
        RECT 114.965 15.355 117.555 16.615 ;
        RECT 115.885 14.265 117.555 16.615 ;
        RECT 115.035 14.555 115.205 16.615 ;
        RECT 114.195 14.555 114.365 15.525 ;
        RECT 114.02 15.355 114.35 16.285 ;
        RECT 113.275 14.555 113.605 15.525 ;
        RECT 113.075 15.355 113.43 15.945 ;
        RECT 112.435 14.555 112.765 15.525 ;
        RECT 111.595 14.555 111.925 15.525 ;
        RECT 110.755 14.205 111.085 15.525 ;
        RECT 109.675 13.725 110.195 17.155 ;
        RECT 108.985 14.265 110.195 16.615 ;
        RECT 108.095 14.205 108.425 16.675 ;
        RECT 107.255 14.555 107.585 16.325 ;
        RECT 106.415 14.555 106.745 16.325 ;
        RECT 105.575 14.555 105.905 16.325 ;
        RECT 104.815 14.555 104.985 16.325 ;
        RECT 103.975 14.555 104.145 16.325 ;
        RECT 103.005 14.19 103.295 16.69 ;
        RECT 102.085 13.745 102.835 17.135 ;
        RECT 101.165 14.265 102.835 16.615 ;
        RECT 101.625 13.745 102.835 16.615 ;
        RECT 100.245 14.265 102.835 15.525 ;
        RECT 99.785 15.355 100.995 17.135 ;
        RECT 96.565 14.265 100.075 15.525 ;
        RECT 98.405 15.355 100.995 16.615 ;
        RECT 98.385 13.745 100.075 15.525 ;
        RECT 96.09 15.355 96.445 15.945 ;
        RECT 95.62 14.595 95.95 15.525 ;
        RECT 95.17 15.355 95.5 16.285 ;
        RECT 94.675 14.935 95.03 15.525 ;
        RECT 94.035 15.355 94.555 17.155 ;
        RECT 93.345 15.355 94.555 16.615 ;
        RECT 92.425 15.355 93.175 17.135 ;
        RECT 91.505 14.265 92.715 16.615 ;
        RECT 92.195 13.725 92.715 16.615 ;
        RECT 90.125 13.745 91.335 17.135 ;
        RECT 88.745 14.265 91.335 16.615 ;
        RECT 88.285 14.19 88.575 16.69 ;
        RECT 87.595 13.725 88.115 17.155 ;
        RECT 86.905 14.265 88.115 16.615 ;
        RECT 85.985 13.745 86.735 17.135 ;
        RECT 85.065 14.265 86.735 16.615 ;
        RECT 79.545 14.265 84.89 15.525 ;
        RECT 82.295 13.745 84.89 15.525 ;
        RECT 82.75 13.745 83.105 15.945 ;
        RECT 81.83 14.265 82.16 16.285 ;
        RECT 80.465 14.265 81.215 17.135 ;
        RECT 79.545 14.265 81.215 16.615 ;
        RECT 74.025 14.265 79.37 15.525 ;
        RECT 76.775 13.745 79.37 15.525 ;
        RECT 78.655 13.745 78.985 16.675 ;
        RECT 77.815 13.745 78.145 16.325 ;
        RECT 76.975 13.745 77.305 16.325 ;
        RECT 76.135 14.265 76.465 16.325 ;
        RECT 75.375 14.265 75.545 16.325 ;
        RECT 74.535 14.265 74.705 16.325 ;
        RECT 73.565 14.19 73.855 16.69 ;
        RECT 72.875 15.355 73.395 17.155 ;
        RECT 72.185 15.355 73.395 16.615 ;
        RECT 71.265 14.265 72.475 15.525 ;
        RECT 71.955 13.725 72.475 15.525 ;
        RECT 70.375 14.205 70.705 15.525 ;
        RECT 69.87 15.355 70.225 15.945 ;
        RECT 69.535 14.555 69.865 15.525 ;
        RECT 68.95 15.355 69.28 16.285 ;
        RECT 68.695 14.555 69.025 15.525 ;
        RECT 67.585 15.355 68.335 17.135 ;
        RECT 67.855 14.555 68.185 17.135 ;
        RECT 66.665 15.355 68.335 16.615 ;
        RECT 67.095 14.555 67.265 16.615 ;
        RECT 66.255 14.555 66.425 15.525 ;
        RECT 65.765 15.355 65.935 16.535 ;
        RECT 64.365 14.265 65.575 15.525 ;
        RECT 65.055 13.725 65.575 15.525 ;
        RECT 64.71 14.265 65.025 16.025 ;
        RECT 62.83 15.355 63 16.325 ;
        RECT 62.05 14.935 62.405 15.525 ;
        RECT 61.13 14.595 61.46 15.525 ;
        RECT 60.66 15.355 60.925 15.985 ;
        RECT 59.305 14.265 60.515 15.525 ;
        RECT 59.995 13.725 60.515 15.525 ;
        RECT 59.735 14.265 60.065 16.025 ;
        RECT 58.845 14.19 59.135 16.69 ;
        RECT 58.155 13.745 58.675 17.155 ;
        RECT 57.465 14.265 58.675 16.615 ;
        RECT 57.925 13.745 58.675 16.615 ;
        RECT 57.005 14.265 58.675 15.525 ;
        RECT 54.245 14.265 56.835 15.525 ;
        RECT 55.625 13.745 56.835 15.525 ;
        RECT 56.565 13.745 56.735 16.535 ;
        RECT 55.51 14.265 55.825 16.025 ;
        RECT 53.63 15.355 53.8 16.325 ;
        RECT 53.3 14.595 53.63 15.525 ;
        RECT 52.355 14.935 52.71 15.525 ;
        RECT 51.46 15.355 51.725 15.985 ;
        RECT 50.535 15.355 50.865 16.025 ;
        RECT 47.805 14.265 50.395 15.525 ;
        RECT 49.185 13.745 50.395 15.525 ;
        RECT 49.185 13.745 49.935 17.135 ;
        RECT 48.265 14.265 49.935 16.615 ;
        RECT 47.32 15.355 47.65 16.285 ;
        RECT 46.865 14.555 47.145 15.525 ;
        RECT 46.375 15.355 46.73 15.945 ;
        RECT 44.125 14.19 44.415 16.69 ;
        RECT 42.745 14.265 43.955 17.135 ;
        RECT 43.435 13.725 43.955 17.135 ;
        RECT 41.365 15.355 43.955 16.615 ;
        RECT 40.905 14.265 42.575 15.525 ;
        RECT 41.825 13.745 42.575 16.615 ;
        RECT 38.145 14.265 40.735 15.525 ;
        RECT 39.525 13.745 40.735 15.525 ;
        RECT 40.515 13.745 40.685 16.325 ;
        RECT 39.675 13.745 39.845 16.325 ;
        RECT 38.755 14.265 39.085 16.325 ;
        RECT 37.915 15.355 38.245 16.325 ;
        RECT 37.295 14.555 37.465 15.525 ;
        RECT 37.075 15.355 37.405 16.325 ;
        RECT 36.455 14.555 36.625 15.525 ;
        RECT 36.235 15.355 36.565 16.675 ;
        RECT 35.535 14.555 35.865 15.525 ;
        RECT 34.695 14.555 35.025 15.525 ;
        RECT 34.495 15.355 34.825 16.675 ;
        RECT 33.855 14.555 34.185 15.525 ;
        RECT 33.655 15.355 33.985 16.325 ;
        RECT 33.015 14.205 33.345 15.525 ;
        RECT 32.815 15.355 33.145 16.325 ;
        RECT 29.865 14.265 32.455 15.525 ;
        RECT 31.245 13.745 32.455 15.525 ;
        RECT 31.975 13.745 32.305 16.325 ;
        RECT 31.215 14.265 31.385 16.325 ;
        RECT 30.375 14.265 30.545 16.325 ;
        RECT 29.405 14.19 29.695 16.69 ;
        RECT 28.485 13.745 29.235 17.135 ;
        RECT 27.565 14.265 29.235 16.615 ;
        RECT 26.185 13.745 27.395 17.135 ;
        RECT 24.805 14.265 27.395 16.615 ;
        RECT 23.915 14.205 24.245 16.675 ;
        RECT 23.075 14.555 23.405 16.325 ;
        RECT 22.235 14.555 22.565 16.325 ;
        RECT 21.395 14.555 21.725 16.325 ;
        RECT 20.635 14.555 20.805 16.325 ;
        RECT 19.795 14.555 19.965 16.325 ;
        RECT 18.595 13.725 19.115 17.155 ;
        RECT 17.905 14.265 19.115 16.615 ;
        RECT 16.525 13.745 17.735 17.135 ;
        RECT 15.145 14.265 17.735 16.615 ;
        RECT 14.685 14.19 14.975 16.69 ;
        RECT 13.995 13.725 14.515 17.155 ;
        RECT 13.305 14.265 14.515 16.615 ;
        RECT 11.925 13.745 13.135 17.135 ;
        RECT 10.545 14.265 13.135 16.615 ;
        RECT 10 20.795 189.86 20.965 ;
        RECT 189.025 19.63 189.315 22.13 ;
        RECT 188.105 19.185 188.855 22.575 ;
        RECT 187.185 19.705 188.855 22.055 ;
        RECT 187.645 19.185 188.855 22.055 ;
        RECT 186.265 19.705 188.855 20.965 ;
        RECT 185.805 20.795 187.015 22.575 ;
        RECT 182.585 19.705 186.095 20.965 ;
        RECT 184.425 20.795 187.015 22.055 ;
        RECT 184.405 19.185 186.095 20.965 ;
        RECT 183.525 19.705 183.695 21.975 ;
        RECT 182.47 20.795 182.785 21.465 ;
        RECT 177.065 19.705 182.41 20.965 ;
        RECT 179.815 19.185 182.41 20.965 ;
        RECT 180.59 19.185 180.76 21.765 ;
        RECT 178.42 19.705 178.685 21.425 ;
        RECT 177.495 19.705 177.825 21.465 ;
        RECT 176.605 19.63 176.895 22.13 ;
        RECT 175.915 19.185 176.435 22.595 ;
        RECT 175.225 19.705 176.435 22.055 ;
        RECT 175.685 19.185 176.435 22.055 ;
        RECT 174.765 19.705 176.435 20.965 ;
        RECT 174.305 20.795 175.055 22.575 ;
        RECT 174.255 20.37 174.59 22.055 ;
        RECT 173.385 20.795 175.055 22.055 ;
        RECT 173.365 20.015 173.695 20.965 ;
        RECT 172.875 20.795 173.21 21.39 ;
        RECT 171.985 20.795 172.315 21.745 ;
        RECT 172.025 19.785 172.195 21.745 ;
        RECT 170.97 20.295 171.285 20.965 ;
        RECT 170.605 20.795 170.935 21.725 ;
        RECT 169.09 19.995 169.26 20.965 ;
        RECT 168.805 20.795 168.975 21.975 ;
        RECT 167.75 20.795 168.065 21.465 ;
        RECT 166.92 20.335 167.185 20.965 ;
        RECT 165.995 20.295 166.325 20.965 ;
        RECT 165.87 20.795 166.04 21.765 ;
        RECT 164.335 20.335 164.66 20.965 ;
        RECT 163.7 20.795 163.965 21.425 ;
        RECT 162.915 20.335 163.185 20.965 ;
        RECT 162.775 20.795 163.105 21.465 ;
        RECT 161.885 19.63 162.175 22.13 ;
        RECT 160.505 19.705 161.715 20.965 ;
        RECT 161.195 19.165 161.715 20.965 ;
        RECT 160.065 20.795 160.235 21.975 ;
        RECT 159.605 19.785 159.775 20.965 ;
        RECT 159.01 20.795 159.325 21.465 ;
        RECT 158.55 20.295 158.865 20.965 ;
        RECT 157.13 20.795 157.3 21.765 ;
        RECT 156.67 19.995 156.84 20.965 ;
        RECT 154.96 20.795 155.225 21.425 ;
        RECT 154.5 20.335 154.765 20.965 ;
        RECT 154.035 20.795 154.365 21.465 ;
        RECT 153.575 20.295 153.905 20.965 ;
        RECT 152.915 20.795 153.435 22.595 ;
        RECT 147.625 19.705 152.97 20.965 ;
        RECT 152.225 20.795 153.435 22.055 ;
        RECT 150.375 19.185 152.97 20.965 ;
        RECT 151.305 19.185 152.055 22.575 ;
        RECT 150.385 19.185 152.055 22.055 ;
        RECT 149.005 19.705 150.215 22.575 ;
        RECT 147.625 19.705 150.215 22.055 ;
        RECT 147.165 19.63 147.455 22.13 ;
        RECT 146.475 20.795 146.995 22.595 ;
        RECT 145.785 20.795 146.995 22.055 ;
        RECT 145.3 20.035 145.63 20.965 ;
        RECT 143.925 20.795 145.615 22.575 ;
        RECT 144.355 20.375 144.71 22.575 ;
        RECT 142.105 20.795 145.615 22.055 ;
        RECT 140.265 19.705 141.475 20.965 ;
        RECT 140.955 19.165 141.475 20.965 ;
        RECT 141.205 19.165 141.375 21.975 ;
        RECT 140.15 20.795 140.465 21.465 ;
        RECT 139.365 19.785 139.535 20.965 ;
        RECT 138.31 20.295 138.625 20.965 ;
        RECT 138.27 20.795 138.44 21.765 ;
        RECT 136.43 19.995 136.6 20.965 ;
        RECT 136.1 20.795 136.365 21.425 ;
        RECT 135.175 20.795 135.505 21.465 ;
        RECT 134.26 20.335 134.525 20.965 ;
        RECT 133.805 20.795 134.135 21.725 ;
        RECT 133.335 20.295 133.665 20.965 ;
        RECT 132.445 19.63 132.735 22.13 ;
        RECT 131.065 19.705 132.275 20.965 ;
        RECT 131.755 19.165 132.275 20.965 ;
        RECT 131.085 19.705 131.255 21.975 ;
        RECT 125.545 19.705 130.89 20.965 ;
        RECT 128.295 19.185 130.89 20.965 ;
        RECT 130.03 19.185 130.345 21.465 ;
        RECT 128.15 19.705 128.32 21.765 ;
        RECT 125.98 19.705 126.245 21.425 ;
        RECT 125.055 20.795 125.385 21.465 ;
        RECT 124.645 19.785 124.815 20.965 ;
        RECT 123.245 20.795 124.455 22.575 ;
        RECT 123.59 20.295 123.905 22.575 ;
        RECT 121.865 20.795 124.455 22.055 ;
        RECT 121.71 19.995 121.88 20.965 ;
        RECT 120.005 20.795 121.695 22.575 ;
        RECT 118.185 20.795 121.695 22.055 ;
        RECT 119.54 20.335 119.805 22.055 ;
        RECT 118.615 20.295 118.945 22.055 ;
        RECT 117.725 19.63 118.015 22.13 ;
        RECT 114.965 19.705 117.555 20.965 ;
        RECT 116.345 19.185 117.555 20.965 ;
        RECT 116.825 19.185 116.995 21.975 ;
        RECT 115.77 19.705 116.085 21.465 ;
        RECT 114.115 19.995 114.285 20.965 ;
        RECT 113.89 20.795 114.06 21.765 ;
        RECT 113.275 19.995 113.445 20.965 ;
        RECT 112.355 19.995 112.685 20.965 ;
        RECT 111.72 20.795 111.985 21.425 ;
        RECT 111.515 19.995 111.845 20.965 ;
        RECT 110.795 20.795 111.125 21.465 ;
        RECT 110.675 19.995 111.005 20.965 ;
        RECT 109.675 20.795 110.195 22.595 ;
        RECT 109.835 19.645 110.165 22.595 ;
        RECT 108.985 20.795 110.195 22.055 ;
        RECT 108.065 19.705 109.275 20.965 ;
        RECT 108.755 19.165 109.275 20.965 ;
        RECT 106.215 20.795 108.81 22.575 ;
        RECT 106.225 19.705 107.895 22.575 ;
        RECT 107.145 19.185 107.895 22.575 ;
        RECT 103.465 20.795 108.81 22.055 ;
        RECT 103.465 19.705 106.055 22.055 ;
        RECT 104.845 19.185 106.055 22.055 ;
        RECT 103.005 19.63 103.295 22.13 ;
        RECT 101.165 19.705 102.835 20.965 ;
        RECT 102.085 19.185 102.835 20.965 ;
        RECT 102.105 19.185 102.275 21.975 ;
        RECT 101.05 20.795 101.365 21.465 ;
        RECT 100.265 19.785 100.435 20.965 ;
        RECT 99.21 20.295 99.525 20.965 ;
        RECT 99.17 20.795 99.34 21.765 ;
        RECT 97.33 19.995 97.5 20.965 ;
        RECT 97 20.795 97.265 21.425 ;
        RECT 96.075 20.795 96.405 21.465 ;
        RECT 94.955 20.795 95.475 22.595 ;
        RECT 95.16 20.335 95.425 22.595 ;
        RECT 94.265 20.795 95.475 22.055 ;
        RECT 94.235 20.295 94.565 20.965 ;
        RECT 91.495 20.795 94.09 22.575 ;
        RECT 92.425 19.705 93.635 22.575 ;
        RECT 93.115 19.165 93.635 22.575 ;
        RECT 88.745 19.705 92.255 22.055 ;
        RECT 90.565 19.185 92.255 22.055 ;
        RECT 88.285 19.63 88.575 22.13 ;
        RECT 86.445 19.705 88.115 20.965 ;
        RECT 87.365 19.185 88.115 20.965 ;
        RECT 87.385 19.185 87.555 21.975 ;
        RECT 86.33 20.795 86.645 21.465 ;
        RECT 85.5 20.035 85.83 20.965 ;
        RECT 84.555 20.375 84.91 20.965 ;
        RECT 84.45 20.795 84.62 21.765 ;
        RECT 82.28 20.795 82.545 21.425 ;
        RECT 81.865 19.785 82.035 20.965 ;
        RECT 81.355 20.795 81.685 21.465 ;
        RECT 80.81 20.295 81.125 20.965 ;
        RECT 79.985 20.795 80.315 21.725 ;
        RECT 76.775 20.795 79.37 22.575 ;
        RECT 78.93 19.995 79.1 22.575 ;
        RECT 76.76 20.335 77.025 22.055 ;
        RECT 74.025 20.795 79.37 22.055 ;
        RECT 75.835 20.295 76.165 22.055 ;
        RECT 74.025 19.705 75.235 22.055 ;
        RECT 74.715 19.165 75.235 22.055 ;
        RECT 73.565 19.63 73.855 22.13 ;
        RECT 72.185 19.705 73.395 20.965 ;
        RECT 72.875 19.165 73.395 20.965 ;
        RECT 72.665 19.705 72.835 21.975 ;
        RECT 71.61 20.795 71.925 21.465 ;
        RECT 69.87 20.375 70.225 20.965 ;
        RECT 69.73 20.795 69.9 21.765 ;
        RECT 68.95 20.035 69.28 20.965 ;
        RECT 66.665 19.705 68.335 20.965 ;
        RECT 67.585 19.185 68.335 20.965 ;
        RECT 67.56 19.705 67.825 21.425 ;
        RECT 66.635 20.795 66.965 21.465 ;
        RECT 65.285 20.795 66.035 22.575 ;
        RECT 65.765 19.785 65.935 22.575 ;
        RECT 64.365 20.795 66.035 22.055 ;
        RECT 64.71 20.295 65.025 22.055 ;
        RECT 62.985 20.795 64.195 22.575 ;
        RECT 62.83 19.995 63 22.055 ;
        RECT 61.605 20.795 64.195 22.055 ;
        RECT 60.665 20.795 60.995 21.725 ;
        RECT 60.66 20.335 60.925 20.965 ;
        RECT 59.735 20.295 60.065 20.965 ;
        RECT 58.845 19.63 59.135 22.13 ;
        RECT 57.005 19.705 58.675 20.965 ;
        RECT 57.925 19.185 58.675 20.965 ;
        RECT 57.945 19.185 58.115 21.975 ;
        RECT 56.89 20.795 57.205 21.465 ;
        RECT 56.105 19.785 56.275 20.965 ;
        RECT 55.05 20.295 55.365 20.965 ;
        RECT 55.01 20.795 55.18 21.765 ;
        RECT 53.17 19.995 53.34 20.965 ;
        RECT 52.84 20.795 53.105 21.425 ;
        RECT 51.915 20.795 52.245 21.465 ;
        RECT 50.565 20.795 51.315 22.575 ;
        RECT 51 20.335 51.265 22.575 ;
        RECT 49.645 20.795 51.315 22.055 ;
        RECT 50.075 20.295 50.405 22.055 ;
        RECT 48.265 19.705 49.475 20.965 ;
        RECT 48.955 19.165 49.475 20.965 ;
        RECT 48.7 19.705 49.03 21.725 ;
        RECT 47.755 20.795 48.11 21.385 ;
        RECT 44.585 19.705 48.095 20.965 ;
        RECT 46.405 19.185 48.095 20.965 ;
        RECT 45.275 19.705 45.795 22.595 ;
        RECT 44.585 19.705 45.795 22.055 ;
        RECT 44.125 19.63 44.415 22.13 ;
        RECT 43.435 19.165 43.955 22.595 ;
        RECT 42.745 19.705 43.955 22.055 ;
        RECT 41.825 19.185 42.575 22.575 ;
        RECT 40.905 19.705 42.575 22.055 ;
        RECT 38.135 19.185 40.73 22.575 ;
        RECT 35.385 19.705 40.73 22.055 ;
        RECT 32.615 19.185 35.21 22.575 ;
        RECT 29.865 19.705 35.21 22.055 ;
        RECT 29.405 19.63 29.695 22.13 ;
        RECT 28.715 19.165 29.235 22.595 ;
        RECT 28.025 19.705 29.235 22.055 ;
        RECT 27.105 19.185 27.855 22.575 ;
        RECT 26.185 19.705 27.855 22.055 ;
        RECT 23.415 19.185 26.01 22.575 ;
        RECT 20.665 19.705 26.01 22.055 ;
        RECT 17.895 19.185 20.49 22.575 ;
        RECT 15.145 19.705 20.49 22.055 ;
        RECT 14.685 19.63 14.975 22.13 ;
        RECT 13.995 19.165 14.515 22.595 ;
        RECT 13.305 19.705 14.515 22.055 ;
        RECT 11.925 19.185 13.135 22.575 ;
        RECT 10.545 19.705 13.135 22.055 ;
        RECT 10 26.235 189.86 26.405 ;
        RECT 189.025 25.07 189.315 27.57 ;
        RECT 187.645 25.145 188.855 28.015 ;
        RECT 188.335 24.605 188.855 28.015 ;
        RECT 186.265 26.235 188.855 27.495 ;
        RECT 185.805 25.145 187.475 26.405 ;
        RECT 186.725 24.625 187.475 27.495 ;
        RECT 184.405 26.235 186.095 28.015 ;
        RECT 184.915 25.085 185.245 28.015 ;
        RECT 184.075 25.435 184.405 27.495 ;
        RECT 182.585 26.235 186.095 27.495 ;
        RECT 183.235 25.435 183.565 27.495 ;
        RECT 182.395 25.435 182.725 26.405 ;
        RECT 179.815 26.235 182.41 28.015 ;
        RECT 181.635 25.435 181.805 28.015 ;
        RECT 180.795 25.435 180.965 28.015 ;
        RECT 178.905 25.145 180.115 27.495 ;
        RECT 179.595 24.605 180.115 27.495 ;
        RECT 177.065 26.235 182.41 27.495 ;
        RECT 177.065 25.145 178.735 27.495 ;
        RECT 177.985 24.625 178.735 27.495 ;
        RECT 176.605 25.07 176.895 27.57 ;
        RECT 175.915 24.625 176.435 28.035 ;
        RECT 175.225 25.145 176.435 27.495 ;
        RECT 175.685 24.625 176.435 27.495 ;
        RECT 174.765 25.145 176.435 26.405 ;
        RECT 174.305 26.235 175.055 28.015 ;
        RECT 172.005 25.145 174.595 26.405 ;
        RECT 173.385 24.625 174.595 27.495 ;
        RECT 170.615 26.235 173.21 28.015 ;
        RECT 171.055 25.525 171.385 28.015 ;
        RECT 167.865 26.235 173.21 27.495 ;
        RECT 169.685 25.505 170.025 27.495 ;
        RECT 167.865 25.145 169.075 27.495 ;
        RECT 168.555 24.605 169.075 27.495 ;
        RECT 165.095 24.625 167.69 28.015 ;
        RECT 162.345 25.145 167.69 27.495 ;
        RECT 161.885 25.07 162.175 27.57 ;
        RECT 161.195 24.605 161.715 28.035 ;
        RECT 160.505 25.145 161.715 27.495 ;
        RECT 158.665 25.145 160.335 26.405 ;
        RECT 159.585 24.625 160.335 26.405 ;
        RECT 159.56 25.145 159.89 27.165 ;
        RECT 158.615 26.235 158.97 26.825 ;
        RECT 156.35 25.815 156.705 26.405 ;
        RECT 154.965 26.235 156.655 28.015 ;
        RECT 155.43 25.475 155.76 28.015 ;
        RECT 153.145 26.235 156.655 27.495 ;
        RECT 153.145 25.145 154.815 27.495 ;
        RECT 154.065 24.625 154.815 27.495 ;
        RECT 150.375 26.235 152.97 28.015 ;
        RECT 152.295 25.435 152.465 28.015 ;
        RECT 151.455 25.435 151.625 28.015 ;
        RECT 150.535 25.435 150.865 28.015 ;
        RECT 147.625 26.235 152.97 27.495 ;
        RECT 149.695 25.435 150.025 27.495 ;
        RECT 148.855 25.435 149.185 27.495 ;
        RECT 148.015 25.085 148.345 27.495 ;
        RECT 147.165 25.07 147.455 27.57 ;
        RECT 146.245 26.235 146.995 28.015 ;
        RECT 141.645 25.145 146.99 26.405 ;
        RECT 145.325 26.235 146.995 27.495 ;
        RECT 144.395 24.625 146.99 26.405 ;
        RECT 143.945 25.145 145.155 28.015 ;
        RECT 142.565 25.145 145.155 27.495 ;
        RECT 141.665 25.145 141.835 27.415 ;
        RECT 140.61 26.235 140.925 26.905 ;
        RECT 139.33 25.815 139.685 26.405 ;
        RECT 138.73 26.235 138.9 27.205 ;
        RECT 138.41 25.475 138.74 26.405 ;
        RECT 136.585 25.145 137.795 26.405 ;
        RECT 137.275 24.605 137.795 26.405 ;
        RECT 136.56 26.235 136.825 26.865 ;
        RECT 132.905 25.145 136.415 26.405 ;
        RECT 134.725 24.625 136.415 26.405 ;
        RECT 135.635 24.625 135.965 26.905 ;
        RECT 133.595 25.145 134.115 28.035 ;
        RECT 132.905 25.145 134.115 27.495 ;
        RECT 132.445 25.07 132.735 27.57 ;
        RECT 131.065 25.145 132.275 26.405 ;
        RECT 131.755 24.605 132.275 26.405 ;
        RECT 131.085 25.145 131.255 27.415 ;
        RECT 125.545 25.145 130.89 26.405 ;
        RECT 128.295 24.625 130.89 26.405 ;
        RECT 130.03 24.625 130.345 26.905 ;
        RECT 128.15 25.145 128.32 27.205 ;
        RECT 125.98 25.145 126.245 26.865 ;
        RECT 125.055 26.235 125.385 26.905 ;
        RECT 124.645 25.225 124.815 26.405 ;
        RECT 123.935 26.235 124.455 28.035 ;
        RECT 123.245 26.235 124.455 27.495 ;
        RECT 123.59 25.735 123.905 27.495 ;
        RECT 122.3 26.235 122.63 27.165 ;
        RECT 121.71 25.435 121.88 26.405 ;
        RECT 121.355 26.235 121.71 26.825 ;
        RECT 119.54 25.775 119.805 26.405 ;
        RECT 118.875 26.235 119.395 28.035 ;
        RECT 118.615 25.735 118.945 27.495 ;
        RECT 118.185 26.235 119.395 27.495 ;
        RECT 117.725 25.07 118.015 27.57 ;
        RECT 117.035 24.605 117.555 28.035 ;
        RECT 116.345 25.145 117.555 27.495 ;
        RECT 115.425 26.235 116.175 28.015 ;
        RECT 115.4 25.475 115.73 27.495 ;
        RECT 114.505 26.235 116.175 27.495 ;
        RECT 114.455 25.815 114.81 26.405 ;
        RECT 111.735 26.235 114.33 28.015 ;
        RECT 108.985 25.145 112.495 27.495 ;
        RECT 110.805 24.625 112.495 27.495 ;
        RECT 106.215 24.625 108.81 28.015 ;
        RECT 103.465 25.145 108.81 27.495 ;
        RECT 103.005 25.07 103.295 27.57 ;
        RECT 102.315 24.625 102.835 28.035 ;
        RECT 101.625 25.145 102.835 27.495 ;
        RECT 102.085 24.625 102.835 27.495 ;
        RECT 101.165 25.145 102.835 26.405 ;
        RECT 100.705 26.235 101.455 28.015 ;
        RECT 98.405 25.145 100.995 26.405 ;
        RECT 99.785 24.625 100.995 27.495 ;
        RECT 97.015 26.235 99.61 28.015 ;
        RECT 97.505 25.225 97.675 28.015 ;
        RECT 94.265 26.235 99.61 27.495 ;
        RECT 96.45 25.735 96.765 27.495 ;
        RECT 94.57 25.435 94.74 27.495 ;
        RECT 91.495 26.235 94.09 28.015 ;
        RECT 92.4 25.775 92.665 28.015 ;
        RECT 91.475 25.735 91.805 27.495 ;
        RECT 88.745 26.235 94.09 27.495 ;
        RECT 88.745 25.145 89.955 27.495 ;
        RECT 89.435 24.605 89.955 27.495 ;
        RECT 88.285 25.07 88.575 27.57 ;
        RECT 87.595 24.625 88.115 28.035 ;
        RECT 86.905 24.625 88.115 27.495 ;
        RECT 84.605 25.145 88.115 26.405 ;
        RECT 86.425 24.625 88.115 26.405 ;
        RECT 85.985 25.145 86.735 28.015 ;
        RECT 85.065 25.145 86.735 27.495 ;
        RECT 82.295 26.235 84.89 28.015 ;
        RECT 83.705 25.225 83.875 28.015 ;
        RECT 82.65 25.735 82.965 28.015 ;
        RECT 79.545 26.235 84.89 27.495 ;
        RECT 80.77 25.435 80.94 27.495 ;
        RECT 76.775 26.235 79.37 28.015 ;
        RECT 78.6 25.775 78.865 28.015 ;
        RECT 77.675 25.735 78.005 28.015 ;
        RECT 75.865 25.145 77.075 27.495 ;
        RECT 76.555 24.605 77.075 27.495 ;
        RECT 74.025 26.235 79.37 27.495 ;
        RECT 74.025 25.145 75.695 27.495 ;
        RECT 74.945 24.625 75.695 27.495 ;
        RECT 73.565 25.07 73.855 27.57 ;
        RECT 72.875 26.235 73.395 28.035 ;
        RECT 72.185 26.235 73.395 27.495 ;
        RECT 71.265 25.145 72.475 26.405 ;
        RECT 71.955 24.605 72.475 26.405 ;
        RECT 70.375 25.085 70.705 26.405 ;
        RECT 69.87 26.235 70.225 26.825 ;
        RECT 69.535 25.435 69.865 26.405 ;
        RECT 68.95 26.235 69.28 27.165 ;
        RECT 68.695 25.435 69.025 26.405 ;
        RECT 67.585 26.235 68.335 28.015 ;
        RECT 67.855 25.435 68.185 28.015 ;
        RECT 66.665 26.235 68.335 27.495 ;
        RECT 67.095 25.435 67.265 27.495 ;
        RECT 66.255 25.435 66.425 26.405 ;
        RECT 65.765 26.235 65.935 27.415 ;
        RECT 62.985 25.145 65.575 26.405 ;
        RECT 64.365 24.625 65.575 26.405 ;
        RECT 64.71 24.625 65.025 26.905 ;
        RECT 62.83 26.235 63 27.205 ;
        RECT 59.305 25.145 62.815 26.405 ;
        RECT 61.125 24.625 62.815 26.405 ;
        RECT 60.66 25.145 60.925 26.865 ;
        RECT 59.735 25.145 60.065 26.905 ;
        RECT 58.845 25.07 59.135 27.57 ;
        RECT 56.985 26.235 58.675 28.015 ;
        RECT 57.925 24.625 58.675 28.015 ;
        RECT 57.005 25.145 58.675 28.015 ;
        RECT 55.165 26.235 58.675 27.495 ;
        RECT 56.105 25.225 56.275 27.495 ;
        RECT 55.05 25.735 55.365 26.405 ;
        RECT 52.395 26.235 54.99 28.015 ;
        RECT 53.17 25.435 53.34 28.015 ;
        RECT 49.645 26.235 54.99 27.495 ;
        RECT 51 25.775 51.265 27.495 ;
        RECT 50.075 25.735 50.405 27.495 ;
        RECT 48.265 25.145 49.475 26.405 ;
        RECT 48.955 24.605 49.475 26.405 ;
        RECT 48.7 25.145 49.03 27.165 ;
        RECT 47.755 26.235 48.11 26.825 ;
        RECT 44.585 25.145 48.095 26.405 ;
        RECT 46.405 24.625 48.095 26.405 ;
        RECT 45.275 25.145 45.795 28.035 ;
        RECT 44.585 25.145 45.795 27.495 ;
        RECT 44.125 25.07 44.415 27.57 ;
        RECT 43.435 24.605 43.955 28.035 ;
        RECT 42.745 25.145 43.955 27.495 ;
        RECT 41.825 24.625 42.575 28.015 ;
        RECT 40.905 25.145 42.575 27.495 ;
        RECT 35.385 25.145 40.73 26.405 ;
        RECT 38.135 24.625 40.73 26.405 ;
        RECT 40.055 24.625 40.225 27.205 ;
        RECT 39.215 24.625 39.385 27.205 ;
        RECT 38.295 24.625 38.625 27.205 ;
        RECT 37.455 25.145 37.785 27.205 ;
        RECT 36.615 25.145 36.945 27.205 ;
        RECT 35.775 25.145 36.105 27.555 ;
        RECT 32.615 24.625 35.21 28.015 ;
        RECT 29.865 25.145 35.21 27.495 ;
        RECT 29.405 25.07 29.695 27.57 ;
        RECT 28.715 24.625 29.235 28.035 ;
        RECT 28.025 24.625 29.235 27.495 ;
        RECT 26.645 25.145 29.235 26.405 ;
        RECT 27.105 25.145 27.855 28.015 ;
        RECT 26.185 26.235 27.855 27.495 ;
        RECT 25.755 25.085 26.085 26.405 ;
        RECT 23.415 26.235 26.01 28.015 ;
        RECT 24.915 25.435 25.245 28.015 ;
        RECT 24.075 25.435 24.405 28.015 ;
        RECT 23.235 25.435 23.565 27.495 ;
        RECT 20.665 26.235 26.01 27.495 ;
        RECT 22.475 25.435 22.645 27.495 ;
        RECT 21.635 25.435 21.805 27.495 ;
        RECT 19.745 25.145 20.955 26.405 ;
        RECT 20.435 24.605 20.955 26.405 ;
        RECT 17.895 26.235 20.49 28.015 ;
        RECT 17.905 25.145 19.575 28.015 ;
        RECT 18.825 24.625 19.575 28.015 ;
        RECT 15.145 26.235 20.49 27.495 ;
        RECT 15.145 25.145 17.735 27.495 ;
        RECT 16.525 24.625 17.735 27.495 ;
        RECT 14.685 25.07 14.975 27.57 ;
        RECT 13.995 24.605 14.515 28.035 ;
        RECT 13.305 25.145 14.515 27.495 ;
        RECT 11.925 24.625 13.135 28.015 ;
        RECT 10.545 25.145 13.135 27.495 ;
        RECT 10 31.675 189.86 31.845 ;
        RECT 189.025 30.51 189.315 33.01 ;
        RECT 187.645 30.065 188.855 33.455 ;
        RECT 186.265 30.585 188.855 32.935 ;
        RECT 184.405 30.065 186.095 33.455 ;
        RECT 182.585 30.585 186.095 32.935 ;
        RECT 179.815 30.065 182.41 33.455 ;
        RECT 177.065 30.585 182.41 32.935 ;
        RECT 176.605 30.51 176.895 33.01 ;
        RECT 175.915 30.045 176.435 33.475 ;
        RECT 175.225 30.585 176.435 32.935 ;
        RECT 174.305 30.065 175.055 33.455 ;
        RECT 173.385 30.585 175.055 32.935 ;
        RECT 170.615 30.065 173.21 33.455 ;
        RECT 167.865 30.585 173.21 32.935 ;
        RECT 165.095 30.065 167.69 33.455 ;
        RECT 162.345 30.585 167.69 32.935 ;
        RECT 161.885 30.51 162.175 33.01 ;
        RECT 161.195 30.045 161.715 33.475 ;
        RECT 160.505 30.585 161.715 32.935 ;
        RECT 159.585 30.065 160.335 33.455 ;
        RECT 158.665 30.585 160.335 32.935 ;
        RECT 155.895 30.065 158.49 33.455 ;
        RECT 153.145 30.585 158.49 32.935 ;
        RECT 150.375 30.065 152.97 33.455 ;
        RECT 147.625 30.585 152.97 32.935 ;
        RECT 147.165 30.51 147.455 33.01 ;
        RECT 146.475 31.675 146.995 33.475 ;
        RECT 141.645 30.585 146.99 31.845 ;
        RECT 145.785 31.675 146.995 32.935 ;
        RECT 144.395 30.065 146.99 31.845 ;
        RECT 144.865 30.065 145.615 33.455 ;
        RECT 143.945 30.585 145.615 32.935 ;
        RECT 141.175 31.675 143.77 33.455 ;
        RECT 138.425 31.675 143.77 32.935 ;
        RECT 139.33 31.255 139.685 32.935 ;
        RECT 138.41 30.915 138.74 31.845 ;
        RECT 135.655 31.675 138.25 33.455 ;
        RECT 136.585 30.585 137.795 33.455 ;
        RECT 137.275 30.045 137.795 33.455 ;
        RECT 132.905 30.585 136.415 32.935 ;
        RECT 134.725 30.065 136.415 32.935 ;
        RECT 132.445 30.51 132.735 33.01 ;
        RECT 131.065 30.065 132.275 33.455 ;
        RECT 129.685 30.585 132.275 32.935 ;
        RECT 130.585 30.065 132.275 32.935 ;
        RECT 128.765 30.585 132.275 31.845 ;
        RECT 127.825 31.675 129.515 33.455 ;
        RECT 123.245 30.585 128.59 31.845 ;
        RECT 126.005 31.675 129.515 32.935 ;
        RECT 125.995 30.065 128.59 31.845 ;
        RECT 123.235 31.675 125.83 33.455 ;
        RECT 120.485 31.675 125.83 32.935 ;
        RECT 122.3 30.915 122.63 32.935 ;
        RECT 121.355 31.255 121.71 32.935 ;
        RECT 120.045 31.675 120.275 32.985 ;
        RECT 118.185 30.585 119.395 31.845 ;
        RECT 118.875 30.045 119.395 31.845 ;
        RECT 119.165 30.045 119.375 32.985 ;
        RECT 117.725 30.51 118.015 33.01 ;
        RECT 117.035 30.045 117.555 33.475 ;
        RECT 116.345 30.585 117.555 32.935 ;
        RECT 115.425 30.065 116.175 33.455 ;
        RECT 114.505 30.585 116.175 32.935 ;
        RECT 111.735 30.065 114.33 33.455 ;
        RECT 108.985 30.585 114.33 32.935 ;
        RECT 106.215 30.065 108.81 33.455 ;
        RECT 103.465 30.585 108.81 32.935 ;
        RECT 103.005 30.51 103.295 33.01 ;
        RECT 102.315 31.675 102.835 33.475 ;
        RECT 97.485 30.585 102.83 31.845 ;
        RECT 101.625 31.675 102.835 32.935 ;
        RECT 100.235 30.065 102.83 31.845 ;
        RECT 100.705 30.065 101.455 33.455 ;
        RECT 99.785 30.585 101.455 32.935 ;
        RECT 97.015 31.675 99.61 33.455 ;
        RECT 94.265 31.675 99.61 32.935 ;
        RECT 96.54 30.915 96.87 32.935 ;
        RECT 95.595 31.255 95.95 32.935 ;
        RECT 91.495 31.675 94.09 33.455 ;
        RECT 92.425 30.585 93.635 33.455 ;
        RECT 93.115 30.045 93.635 33.455 ;
        RECT 88.745 30.585 92.255 32.935 ;
        RECT 90.565 30.065 92.255 32.935 ;
        RECT 88.285 30.51 88.575 33.01 ;
        RECT 87.595 30.045 88.115 33.475 ;
        RECT 86.905 30.585 88.115 32.935 ;
        RECT 85.985 30.065 86.735 33.455 ;
        RECT 85.065 30.585 86.735 32.935 ;
        RECT 85.525 30.065 86.735 32.935 ;
        RECT 84.145 30.585 86.735 31.845 ;
        RECT 82.295 31.675 84.89 33.455 ;
        RECT 83.2 30.915 83.53 33.455 ;
        RECT 82.255 31.255 82.61 32.935 ;
        RECT 79.545 31.675 84.89 32.935 ;
        RECT 77.705 30.585 80.295 31.845 ;
        RECT 79.085 30.065 80.295 31.845 ;
        RECT 76.775 31.675 79.37 33.455 ;
        RECT 76.76 30.915 77.09 32.935 ;
        RECT 74.025 31.675 79.37 32.935 ;
        RECT 75.815 31.255 76.17 32.935 ;
        RECT 73.565 30.51 73.855 33.01 ;
        RECT 72.875 30.045 73.395 33.475 ;
        RECT 72.185 30.585 73.395 32.935 ;
        RECT 71.265 31.675 72.015 33.455 ;
        RECT 66.665 30.585 72.01 31.845 ;
        RECT 70.345 31.675 72.015 32.935 ;
        RECT 69.415 30.065 72.01 31.845 ;
        RECT 67.575 30.585 70.17 33.455 ;
        RECT 64.825 31.675 70.17 32.935 ;
        RECT 65.765 30.665 65.935 32.935 ;
        RECT 64.71 31.175 65.025 31.845 ;
        RECT 62.055 31.675 64.65 33.455 ;
        RECT 62.83 30.875 63 33.455 ;
        RECT 59.305 31.675 64.65 32.935 ;
        RECT 60.66 31.215 60.925 32.935 ;
        RECT 59.735 31.175 60.065 32.935 ;
        RECT 58.845 30.51 59.135 33.01 ;
        RECT 57.465 30.065 58.675 33.455 ;
        RECT 56.085 30.585 58.675 32.935 ;
      LAYER met1 ;
        RECT 10 9.76 190 10.24 ;
        RECT 10 15.2 190 15.68 ;
        RECT 10 20.64 190 21.12 ;
        RECT 10 26.08 190 26.56 ;
        RECT 10 31.52 190 32 ;
        RECT 10 36.96 190 37.44 ;
        RECT 10 42.4 190 42.88 ;
        RECT 10 47.84 190 48.32 ;
        RECT 10 53.28 190 53.76 ;
        RECT 10 58.72 190 59.2 ;
      LAYER met4 ;
        RECT 184.55 44.7 185.97 46.7 ;
        RECT 184.55 24.3 185.97 26.3 ;
        RECT 184.79 10 185.73 60 ;
        RECT 179.03 44.7 180.45 46.7 ;
        RECT 179.03 24.3 180.45 26.3 ;
        RECT 179.27 10 180.21 60 ;
        RECT 173.51 44.7 174.93 46.7 ;
        RECT 173.51 24.3 174.93 26.3 ;
        RECT 173.75 10 174.69 60 ;
        RECT 167.99 44.7 169.41 46.7 ;
        RECT 167.99 24.3 169.41 26.3 ;
        RECT 168.23 10 169.17 60 ;
        RECT 162.47 44.7 163.89 46.7 ;
        RECT 162.47 24.3 163.89 26.3 ;
        RECT 162.71 10 163.65 60 ;
        RECT 156.95 44.7 158.37 46.7 ;
        RECT 156.95 24.3 158.37 26.3 ;
        RECT 157.19 10 158.13 60 ;
        RECT 151.43 44.7 152.85 46.7 ;
        RECT 151.43 24.3 152.85 26.3 ;
        RECT 151.67 10 152.61 60 ;
        RECT 145.91 44.7 147.33 46.7 ;
        RECT 145.91 24.3 147.33 26.3 ;
        RECT 146.15 10 147.09 60 ;
        RECT 140.39 44.7 141.81 46.7 ;
        RECT 140.39 24.3 141.81 26.3 ;
        RECT 140.63 10 141.57 60 ;
        RECT 134.87 44.7 136.29 46.7 ;
        RECT 134.87 24.3 136.29 26.3 ;
        RECT 135.11 10 136.05 60 ;
        RECT 129.35 44.7 130.77 46.7 ;
        RECT 129.35 24.3 130.77 26.3 ;
        RECT 129.59 10 130.53 60 ;
        RECT 123.83 44.7 125.25 46.7 ;
        RECT 123.83 24.3 125.25 26.3 ;
        RECT 124.07 10 125.01 60 ;
        RECT 118.31 44.7 119.73 46.7 ;
        RECT 118.31 24.3 119.73 26.3 ;
        RECT 118.55 10 119.49 60 ;
        RECT 112.79 44.7 114.21 46.7 ;
        RECT 112.79 24.3 114.21 26.3 ;
        RECT 113.03 10 113.97 60 ;
        RECT 107.27 44.7 108.69 46.7 ;
        RECT 107.27 24.3 108.69 26.3 ;
        RECT 107.51 10 108.45 60 ;
        RECT 101.75 44.7 103.17 46.7 ;
        RECT 101.75 24.3 103.17 26.3 ;
        RECT 101.99 10 102.93 60 ;
        RECT 96.23 44.7 97.65 46.7 ;
        RECT 96.23 24.3 97.65 26.3 ;
        RECT 96.47 10 97.41 60 ;
        RECT 90.71 44.7 92.13 46.7 ;
        RECT 90.71 24.3 92.13 26.3 ;
        RECT 90.95 10 91.89 60 ;
        RECT 85.19 44.7 86.61 46.7 ;
        RECT 85.19 24.3 86.61 26.3 ;
        RECT 85.43 10 86.37 60 ;
        RECT 79.67 44.7 81.09 46.7 ;
        RECT 79.67 24.3 81.09 26.3 ;
        RECT 79.91 10 80.85 60 ;
        RECT 74.15 44.7 75.57 46.7 ;
        RECT 74.15 24.3 75.57 26.3 ;
        RECT 74.39 10 75.33 60 ;
        RECT 68.63 44.7 70.05 46.7 ;
        RECT 68.63 24.3 70.05 26.3 ;
        RECT 68.87 10 69.81 60 ;
        RECT 63.11 44.7 64.53 46.7 ;
        RECT 63.11 24.3 64.53 26.3 ;
        RECT 63.35 10 64.29 60 ;
        RECT 57.59 44.7 59.01 46.7 ;
        RECT 57.59 24.3 59.01 26.3 ;
        RECT 57.83 10 58.77 60 ;
        RECT 52.07 44.7 53.49 46.7 ;
        RECT 52.07 24.3 53.49 26.3 ;
        RECT 52.31 10 53.25 60 ;
        RECT 46.55 44.7 47.97 46.7 ;
        RECT 46.55 24.3 47.97 26.3 ;
        RECT 46.79 10 47.73 60 ;
        RECT 41.03 44.7 42.45 46.7 ;
        RECT 41.03 24.3 42.45 26.3 ;
        RECT 41.27 10 42.21 60 ;
        RECT 35.51 44.7 36.93 46.7 ;
        RECT 35.51 24.3 36.93 26.3 ;
        RECT 35.75 10 36.69 60 ;
        RECT 29.99 44.7 31.41 46.7 ;
        RECT 29.99 24.3 31.41 26.3 ;
        RECT 30.23 10 31.17 60 ;
        RECT 24.47 44.7 25.89 46.7 ;
        RECT 24.47 24.3 25.89 26.3 ;
        RECT 24.71 10 25.65 60 ;
        RECT 18.95 44.7 20.37 46.7 ;
        RECT 18.95 24.3 20.37 26.3 ;
        RECT 19.19 10 20.13 60 ;
        RECT 13.43 44.7 14.85 46.7 ;
        RECT 13.43 24.3 14.85 26.3 ;
        RECT 13.67 10 14.61 60 ;
      LAYER met3 ;
        RECT 10 12.83 190 13.29 ;
        RECT 10 16.91 190 17.37 ;
        RECT 10 20.99 190 21.45 ;
        RECT 10 25.07 190 25.53 ;
        RECT 10 29.15 190 29.61 ;
        RECT 10 33.23 190 33.69 ;
        RECT 10 37.31 190 37.77 ;
        RECT 10 41.39 190 41.85 ;
        RECT 10 45.47 190 45.93 ;
        RECT 10 49.55 190 50.01 ;
        RECT 10 53.63 190 54.09 ;
        RECT 10 57.71 190 58.17 ;
      LAYER met2 ;
        RECT 188.46 9.98 188.96 60 ;
        RECT 185.7 9.98 186.2 60 ;
        RECT 182.94 9.98 183.44 60 ;
        RECT 180.18 9.98 180.68 60 ;
        RECT 177.42 9.98 177.92 60 ;
        RECT 174.66 9.98 175.16 60 ;
        RECT 171.9 9.98 172.4 60 ;
        RECT 169.14 9.98 169.64 60 ;
        RECT 166.38 9.98 166.88 60 ;
        RECT 163.62 9.98 164.12 60 ;
        RECT 160.86 9.98 161.36 60 ;
        RECT 158.1 9.98 158.6 60 ;
        RECT 155.34 9.98 155.84 60 ;
        RECT 152.58 9.98 153.08 60 ;
        RECT 149.82 9.98 150.32 60 ;
        RECT 147.06 9.98 147.56 60 ;
        RECT 144.3 9.98 144.8 60 ;
        RECT 141.54 9.98 142.04 60 ;
        RECT 138.78 9.98 139.28 60 ;
        RECT 136.02 9.98 136.52 60 ;
        RECT 133.26 9.98 133.76 60 ;
        RECT 130.5 9.98 131 60 ;
        RECT 127.74 9.98 128.24 60 ;
        RECT 124.98 9.98 125.48 60 ;
        RECT 122.22 9.98 122.72 60 ;
        RECT 119.46 9.98 119.96 60 ;
        RECT 116.7 9.98 117.2 60 ;
        RECT 113.94 9.98 114.44 60 ;
        RECT 111.18 9.98 111.68 60 ;
        RECT 108.42 9.98 108.92 60 ;
        RECT 105.66 9.98 106.16 60 ;
        RECT 102.9 9.98 103.4 60 ;
        RECT 100.14 9.98 100.64 60 ;
        RECT 97.38 9.98 97.88 60 ;
        RECT 94.62 9.98 95.12 60 ;
        RECT 91.86 9.98 92.36 60 ;
        RECT 89.1 9.98 89.6 60 ;
        RECT 86.34 9.98 86.84 60 ;
        RECT 83.58 9.98 84.08 60 ;
        RECT 80.82 9.98 81.32 60 ;
        RECT 78.06 9.98 78.56 60 ;
        RECT 75.3 9.98 75.8 60 ;
        RECT 72.54 9.98 73.04 60 ;
        RECT 69.78 9.98 70.28 60 ;
        RECT 67.02 9.98 67.52 60 ;
        RECT 64.26 9.98 64.76 60 ;
        RECT 61.5 9.98 62 60 ;
        RECT 58.74 9.98 59.24 60 ;
        RECT 55.98 9.98 56.48 60 ;
        RECT 53.22 9.98 53.72 60 ;
        RECT 50.46 9.98 50.96 60 ;
        RECT 47.7 9.98 48.2 60 ;
        RECT 44.94 9.98 45.44 60 ;
        RECT 42.18 9.98 42.68 60 ;
        RECT 39.42 9.98 39.92 60 ;
        RECT 36.66 9.98 37.16 60 ;
        RECT 33.9 9.98 34.4 60 ;
        RECT 31.14 9.98 31.64 60 ;
        RECT 28.38 9.98 28.88 60 ;
        RECT 25.62 9.98 26.12 60 ;
        RECT 22.86 9.98 23.36 60 ;
        RECT 20.1 9.98 20.6 60 ;
        RECT 17.34 9.98 17.84 60 ;
        RECT 14.58 9.98 15.08 60 ;
        RECT 11.82 9.98 12.32 60 ;
      LAYER via3 ;
        RECT 13.84 57.84 14.04 58.04 ;
        RECT 13.84 53.76 14.04 53.96 ;
        RECT 13.84 49.68 14.04 49.88 ;
        RECT 13.84 45.6 14.04 45.8 ;
        RECT 13.84 41.52 14.04 41.72 ;
        RECT 13.84 37.44 14.04 37.64 ;
        RECT 13.84 33.36 14.04 33.56 ;
        RECT 13.84 29.28 14.04 29.48 ;
        RECT 13.84 25.2 14.04 25.4 ;
        RECT 13.84 21.12 14.04 21.32 ;
        RECT 13.84 17.04 14.04 17.24 ;
        RECT 13.84 12.96 14.04 13.16 ;
        RECT 14.24 57.84 14.44 58.04 ;
        RECT 14.24 53.76 14.44 53.96 ;
        RECT 14.24 49.68 14.44 49.88 ;
        RECT 14.24 45.6 14.44 45.8 ;
        RECT 14.24 41.52 14.44 41.72 ;
        RECT 14.24 37.44 14.44 37.64 ;
        RECT 14.24 33.36 14.44 33.56 ;
        RECT 14.24 29.28 14.44 29.48 ;
        RECT 14.24 25.2 14.44 25.4 ;
        RECT 14.24 21.12 14.44 21.32 ;
        RECT 14.24 17.04 14.44 17.24 ;
        RECT 14.24 12.96 14.44 13.16 ;
        RECT 19.36 57.84 19.56 58.04 ;
        RECT 19.36 53.76 19.56 53.96 ;
        RECT 19.36 49.68 19.56 49.88 ;
        RECT 19.36 45.6 19.56 45.8 ;
        RECT 19.36 41.52 19.56 41.72 ;
        RECT 19.36 37.44 19.56 37.64 ;
        RECT 19.36 33.36 19.56 33.56 ;
        RECT 19.36 29.28 19.56 29.48 ;
        RECT 19.36 25.2 19.56 25.4 ;
        RECT 19.36 21.12 19.56 21.32 ;
        RECT 19.36 17.04 19.56 17.24 ;
        RECT 19.36 12.96 19.56 13.16 ;
        RECT 19.76 57.84 19.96 58.04 ;
        RECT 19.76 53.76 19.96 53.96 ;
        RECT 19.76 49.68 19.96 49.88 ;
        RECT 19.76 45.6 19.96 45.8 ;
        RECT 19.76 41.52 19.96 41.72 ;
        RECT 19.76 37.44 19.96 37.64 ;
        RECT 19.76 33.36 19.96 33.56 ;
        RECT 19.76 29.28 19.96 29.48 ;
        RECT 19.76 25.2 19.96 25.4 ;
        RECT 19.76 21.12 19.96 21.32 ;
        RECT 19.76 17.04 19.96 17.24 ;
        RECT 19.76 12.96 19.96 13.16 ;
        RECT 24.88 57.84 25.08 58.04 ;
        RECT 24.88 53.76 25.08 53.96 ;
        RECT 24.88 49.68 25.08 49.88 ;
        RECT 24.88 45.6 25.08 45.8 ;
        RECT 24.88 41.52 25.08 41.72 ;
        RECT 24.88 37.44 25.08 37.64 ;
        RECT 24.88 33.36 25.08 33.56 ;
        RECT 24.88 29.28 25.08 29.48 ;
        RECT 24.88 25.2 25.08 25.4 ;
        RECT 24.88 21.12 25.08 21.32 ;
        RECT 24.88 17.04 25.08 17.24 ;
        RECT 24.88 12.96 25.08 13.16 ;
        RECT 25.28 57.84 25.48 58.04 ;
        RECT 25.28 53.76 25.48 53.96 ;
        RECT 25.28 49.68 25.48 49.88 ;
        RECT 25.28 45.6 25.48 45.8 ;
        RECT 25.28 41.52 25.48 41.72 ;
        RECT 25.28 37.44 25.48 37.64 ;
        RECT 25.28 33.36 25.48 33.56 ;
        RECT 25.28 29.28 25.48 29.48 ;
        RECT 25.28 25.2 25.48 25.4 ;
        RECT 25.28 21.12 25.48 21.32 ;
        RECT 25.28 17.04 25.48 17.24 ;
        RECT 25.28 12.96 25.48 13.16 ;
        RECT 30.4 57.84 30.6 58.04 ;
        RECT 30.4 53.76 30.6 53.96 ;
        RECT 30.4 49.68 30.6 49.88 ;
        RECT 30.4 45.6 30.6 45.8 ;
        RECT 30.4 41.52 30.6 41.72 ;
        RECT 30.4 37.44 30.6 37.64 ;
        RECT 30.4 33.36 30.6 33.56 ;
        RECT 30.4 29.28 30.6 29.48 ;
        RECT 30.4 25.2 30.6 25.4 ;
        RECT 30.4 21.12 30.6 21.32 ;
        RECT 30.4 17.04 30.6 17.24 ;
        RECT 30.4 12.96 30.6 13.16 ;
        RECT 30.8 57.84 31 58.04 ;
        RECT 30.8 53.76 31 53.96 ;
        RECT 30.8 49.68 31 49.88 ;
        RECT 30.8 45.6 31 45.8 ;
        RECT 30.8 41.52 31 41.72 ;
        RECT 30.8 37.44 31 37.64 ;
        RECT 30.8 33.36 31 33.56 ;
        RECT 30.8 29.28 31 29.48 ;
        RECT 30.8 25.2 31 25.4 ;
        RECT 30.8 21.12 31 21.32 ;
        RECT 30.8 17.04 31 17.24 ;
        RECT 30.8 12.96 31 13.16 ;
        RECT 35.92 57.84 36.12 58.04 ;
        RECT 35.92 53.76 36.12 53.96 ;
        RECT 35.92 49.68 36.12 49.88 ;
        RECT 35.92 45.6 36.12 45.8 ;
        RECT 35.92 41.52 36.12 41.72 ;
        RECT 35.92 37.44 36.12 37.64 ;
        RECT 35.92 33.36 36.12 33.56 ;
        RECT 35.92 29.28 36.12 29.48 ;
        RECT 35.92 25.2 36.12 25.4 ;
        RECT 35.92 21.12 36.12 21.32 ;
        RECT 35.92 17.04 36.12 17.24 ;
        RECT 35.92 12.96 36.12 13.16 ;
        RECT 36.32 57.84 36.52 58.04 ;
        RECT 36.32 53.76 36.52 53.96 ;
        RECT 36.32 49.68 36.52 49.88 ;
        RECT 36.32 45.6 36.52 45.8 ;
        RECT 36.32 41.52 36.52 41.72 ;
        RECT 36.32 37.44 36.52 37.64 ;
        RECT 36.32 33.36 36.52 33.56 ;
        RECT 36.32 29.28 36.52 29.48 ;
        RECT 36.32 25.2 36.52 25.4 ;
        RECT 36.32 21.12 36.52 21.32 ;
        RECT 36.32 17.04 36.52 17.24 ;
        RECT 36.32 12.96 36.52 13.16 ;
        RECT 41.44 57.84 41.64 58.04 ;
        RECT 41.44 53.76 41.64 53.96 ;
        RECT 41.44 49.68 41.64 49.88 ;
        RECT 41.44 45.6 41.64 45.8 ;
        RECT 41.44 41.52 41.64 41.72 ;
        RECT 41.44 37.44 41.64 37.64 ;
        RECT 41.44 33.36 41.64 33.56 ;
        RECT 41.44 29.28 41.64 29.48 ;
        RECT 41.44 25.2 41.64 25.4 ;
        RECT 41.44 21.12 41.64 21.32 ;
        RECT 41.44 17.04 41.64 17.24 ;
        RECT 41.44 12.96 41.64 13.16 ;
        RECT 41.84 57.84 42.04 58.04 ;
        RECT 41.84 53.76 42.04 53.96 ;
        RECT 41.84 49.68 42.04 49.88 ;
        RECT 41.84 45.6 42.04 45.8 ;
        RECT 41.84 41.52 42.04 41.72 ;
        RECT 41.84 37.44 42.04 37.64 ;
        RECT 41.84 33.36 42.04 33.56 ;
        RECT 41.84 29.28 42.04 29.48 ;
        RECT 41.84 25.2 42.04 25.4 ;
        RECT 41.84 21.12 42.04 21.32 ;
        RECT 41.84 17.04 42.04 17.24 ;
        RECT 41.84 12.96 42.04 13.16 ;
        RECT 46.96 57.84 47.16 58.04 ;
        RECT 46.96 53.76 47.16 53.96 ;
        RECT 46.96 49.68 47.16 49.88 ;
        RECT 46.96 45.6 47.16 45.8 ;
        RECT 46.96 41.52 47.16 41.72 ;
        RECT 46.96 37.44 47.16 37.64 ;
        RECT 46.96 33.36 47.16 33.56 ;
        RECT 46.96 29.28 47.16 29.48 ;
        RECT 46.96 25.2 47.16 25.4 ;
        RECT 46.96 21.12 47.16 21.32 ;
        RECT 46.96 17.04 47.16 17.24 ;
        RECT 46.96 12.96 47.16 13.16 ;
        RECT 47.36 57.84 47.56 58.04 ;
        RECT 47.36 53.76 47.56 53.96 ;
        RECT 47.36 49.68 47.56 49.88 ;
        RECT 47.36 45.6 47.56 45.8 ;
        RECT 47.36 41.52 47.56 41.72 ;
        RECT 47.36 37.44 47.56 37.64 ;
        RECT 47.36 33.36 47.56 33.56 ;
        RECT 47.36 29.28 47.56 29.48 ;
        RECT 47.36 25.2 47.56 25.4 ;
        RECT 47.36 21.12 47.56 21.32 ;
        RECT 47.36 17.04 47.56 17.24 ;
        RECT 47.36 12.96 47.56 13.16 ;
        RECT 52.48 57.84 52.68 58.04 ;
        RECT 52.48 53.76 52.68 53.96 ;
        RECT 52.48 49.68 52.68 49.88 ;
        RECT 52.48 45.6 52.68 45.8 ;
        RECT 52.48 41.52 52.68 41.72 ;
        RECT 52.48 37.44 52.68 37.64 ;
        RECT 52.48 33.36 52.68 33.56 ;
        RECT 52.48 29.28 52.68 29.48 ;
        RECT 52.48 25.2 52.68 25.4 ;
        RECT 52.48 21.12 52.68 21.32 ;
        RECT 52.48 17.04 52.68 17.24 ;
        RECT 52.48 12.96 52.68 13.16 ;
        RECT 52.88 57.84 53.08 58.04 ;
        RECT 52.88 53.76 53.08 53.96 ;
        RECT 52.88 49.68 53.08 49.88 ;
        RECT 52.88 45.6 53.08 45.8 ;
        RECT 52.88 41.52 53.08 41.72 ;
        RECT 52.88 37.44 53.08 37.64 ;
        RECT 52.88 33.36 53.08 33.56 ;
        RECT 52.88 29.28 53.08 29.48 ;
        RECT 52.88 25.2 53.08 25.4 ;
        RECT 52.88 21.12 53.08 21.32 ;
        RECT 52.88 17.04 53.08 17.24 ;
        RECT 52.88 12.96 53.08 13.16 ;
        RECT 58 57.84 58.2 58.04 ;
        RECT 58 53.76 58.2 53.96 ;
        RECT 58 49.68 58.2 49.88 ;
        RECT 58 45.6 58.2 45.8 ;
        RECT 58 41.52 58.2 41.72 ;
        RECT 58 37.44 58.2 37.64 ;
        RECT 58 33.36 58.2 33.56 ;
        RECT 58 29.28 58.2 29.48 ;
        RECT 58 25.2 58.2 25.4 ;
        RECT 58 21.12 58.2 21.32 ;
        RECT 58 17.04 58.2 17.24 ;
        RECT 58 12.96 58.2 13.16 ;
        RECT 58.4 57.84 58.6 58.04 ;
        RECT 58.4 53.76 58.6 53.96 ;
        RECT 58.4 49.68 58.6 49.88 ;
        RECT 58.4 45.6 58.6 45.8 ;
        RECT 58.4 41.52 58.6 41.72 ;
        RECT 58.4 37.44 58.6 37.64 ;
        RECT 58.4 33.36 58.6 33.56 ;
        RECT 58.4 29.28 58.6 29.48 ;
        RECT 58.4 25.2 58.6 25.4 ;
        RECT 58.4 21.12 58.6 21.32 ;
        RECT 58.4 17.04 58.6 17.24 ;
        RECT 58.4 12.96 58.6 13.16 ;
        RECT 63.52 57.84 63.72 58.04 ;
        RECT 63.52 53.76 63.72 53.96 ;
        RECT 63.52 49.68 63.72 49.88 ;
        RECT 63.52 45.6 63.72 45.8 ;
        RECT 63.52 41.52 63.72 41.72 ;
        RECT 63.52 37.44 63.72 37.64 ;
        RECT 63.52 33.36 63.72 33.56 ;
        RECT 63.52 29.28 63.72 29.48 ;
        RECT 63.52 25.2 63.72 25.4 ;
        RECT 63.52 21.12 63.72 21.32 ;
        RECT 63.52 17.04 63.72 17.24 ;
        RECT 63.52 12.96 63.72 13.16 ;
        RECT 63.92 57.84 64.12 58.04 ;
        RECT 63.92 53.76 64.12 53.96 ;
        RECT 63.92 49.68 64.12 49.88 ;
        RECT 63.92 45.6 64.12 45.8 ;
        RECT 63.92 41.52 64.12 41.72 ;
        RECT 63.92 37.44 64.12 37.64 ;
        RECT 63.92 33.36 64.12 33.56 ;
        RECT 63.92 29.28 64.12 29.48 ;
        RECT 63.92 25.2 64.12 25.4 ;
        RECT 63.92 21.12 64.12 21.32 ;
        RECT 63.92 17.04 64.12 17.24 ;
        RECT 63.92 12.96 64.12 13.16 ;
        RECT 69.04 57.84 69.24 58.04 ;
        RECT 69.04 53.76 69.24 53.96 ;
        RECT 69.04 49.68 69.24 49.88 ;
        RECT 69.04 45.6 69.24 45.8 ;
        RECT 69.04 41.52 69.24 41.72 ;
        RECT 69.04 37.44 69.24 37.64 ;
        RECT 69.04 33.36 69.24 33.56 ;
        RECT 69.04 29.28 69.24 29.48 ;
        RECT 69.04 25.2 69.24 25.4 ;
        RECT 69.04 21.12 69.24 21.32 ;
        RECT 69.04 17.04 69.24 17.24 ;
        RECT 69.04 12.96 69.24 13.16 ;
        RECT 69.44 57.84 69.64 58.04 ;
        RECT 69.44 53.76 69.64 53.96 ;
        RECT 69.44 49.68 69.64 49.88 ;
        RECT 69.44 45.6 69.64 45.8 ;
        RECT 69.44 41.52 69.64 41.72 ;
        RECT 69.44 37.44 69.64 37.64 ;
        RECT 69.44 33.36 69.64 33.56 ;
        RECT 69.44 29.28 69.64 29.48 ;
        RECT 69.44 25.2 69.64 25.4 ;
        RECT 69.44 21.12 69.64 21.32 ;
        RECT 69.44 17.04 69.64 17.24 ;
        RECT 69.44 12.96 69.64 13.16 ;
        RECT 74.56 57.84 74.76 58.04 ;
        RECT 74.56 53.76 74.76 53.96 ;
        RECT 74.56 49.68 74.76 49.88 ;
        RECT 74.56 45.6 74.76 45.8 ;
        RECT 74.56 41.52 74.76 41.72 ;
        RECT 74.56 37.44 74.76 37.64 ;
        RECT 74.56 33.36 74.76 33.56 ;
        RECT 74.56 29.28 74.76 29.48 ;
        RECT 74.56 25.2 74.76 25.4 ;
        RECT 74.56 21.12 74.76 21.32 ;
        RECT 74.56 17.04 74.76 17.24 ;
        RECT 74.56 12.96 74.76 13.16 ;
        RECT 74.96 57.84 75.16 58.04 ;
        RECT 74.96 53.76 75.16 53.96 ;
        RECT 74.96 49.68 75.16 49.88 ;
        RECT 74.96 45.6 75.16 45.8 ;
        RECT 74.96 41.52 75.16 41.72 ;
        RECT 74.96 37.44 75.16 37.64 ;
        RECT 74.96 33.36 75.16 33.56 ;
        RECT 74.96 29.28 75.16 29.48 ;
        RECT 74.96 25.2 75.16 25.4 ;
        RECT 74.96 21.12 75.16 21.32 ;
        RECT 74.96 17.04 75.16 17.24 ;
        RECT 74.96 12.96 75.16 13.16 ;
        RECT 80.08 57.84 80.28 58.04 ;
        RECT 80.08 53.76 80.28 53.96 ;
        RECT 80.08 49.68 80.28 49.88 ;
        RECT 80.08 45.6 80.28 45.8 ;
        RECT 80.08 41.52 80.28 41.72 ;
        RECT 80.08 37.44 80.28 37.64 ;
        RECT 80.08 33.36 80.28 33.56 ;
        RECT 80.08 29.28 80.28 29.48 ;
        RECT 80.08 25.2 80.28 25.4 ;
        RECT 80.08 21.12 80.28 21.32 ;
        RECT 80.08 17.04 80.28 17.24 ;
        RECT 80.08 12.96 80.28 13.16 ;
        RECT 80.48 57.84 80.68 58.04 ;
        RECT 80.48 53.76 80.68 53.96 ;
        RECT 80.48 49.68 80.68 49.88 ;
        RECT 80.48 45.6 80.68 45.8 ;
        RECT 80.48 41.52 80.68 41.72 ;
        RECT 80.48 37.44 80.68 37.64 ;
        RECT 80.48 33.36 80.68 33.56 ;
        RECT 80.48 29.28 80.68 29.48 ;
        RECT 80.48 25.2 80.68 25.4 ;
        RECT 80.48 21.12 80.68 21.32 ;
        RECT 80.48 17.04 80.68 17.24 ;
        RECT 80.48 12.96 80.68 13.16 ;
        RECT 85.6 57.84 85.8 58.04 ;
        RECT 85.6 53.76 85.8 53.96 ;
        RECT 85.6 49.68 85.8 49.88 ;
        RECT 85.6 45.6 85.8 45.8 ;
        RECT 85.6 41.52 85.8 41.72 ;
        RECT 85.6 37.44 85.8 37.64 ;
        RECT 85.6 33.36 85.8 33.56 ;
        RECT 85.6 29.28 85.8 29.48 ;
        RECT 85.6 25.2 85.8 25.4 ;
        RECT 85.6 21.12 85.8 21.32 ;
        RECT 85.6 17.04 85.8 17.24 ;
        RECT 85.6 12.96 85.8 13.16 ;
        RECT 86 57.84 86.2 58.04 ;
        RECT 86 53.76 86.2 53.96 ;
        RECT 86 49.68 86.2 49.88 ;
        RECT 86 45.6 86.2 45.8 ;
        RECT 86 41.52 86.2 41.72 ;
        RECT 86 37.44 86.2 37.64 ;
        RECT 86 33.36 86.2 33.56 ;
        RECT 86 29.28 86.2 29.48 ;
        RECT 86 25.2 86.2 25.4 ;
        RECT 86 21.12 86.2 21.32 ;
        RECT 86 17.04 86.2 17.24 ;
        RECT 86 12.96 86.2 13.16 ;
        RECT 91.12 57.84 91.32 58.04 ;
        RECT 91.12 53.76 91.32 53.96 ;
        RECT 91.12 49.68 91.32 49.88 ;
        RECT 91.12 45.6 91.32 45.8 ;
        RECT 91.12 41.52 91.32 41.72 ;
        RECT 91.12 37.44 91.32 37.64 ;
        RECT 91.12 33.36 91.32 33.56 ;
        RECT 91.12 29.28 91.32 29.48 ;
        RECT 91.12 25.2 91.32 25.4 ;
        RECT 91.12 21.12 91.32 21.32 ;
        RECT 91.12 17.04 91.32 17.24 ;
        RECT 91.12 12.96 91.32 13.16 ;
        RECT 91.52 57.84 91.72 58.04 ;
        RECT 91.52 53.76 91.72 53.96 ;
        RECT 91.52 49.68 91.72 49.88 ;
        RECT 91.52 45.6 91.72 45.8 ;
        RECT 91.52 41.52 91.72 41.72 ;
        RECT 91.52 37.44 91.72 37.64 ;
        RECT 91.52 33.36 91.72 33.56 ;
        RECT 91.52 29.28 91.72 29.48 ;
        RECT 91.52 25.2 91.72 25.4 ;
        RECT 91.52 21.12 91.72 21.32 ;
        RECT 91.52 17.04 91.72 17.24 ;
        RECT 91.52 12.96 91.72 13.16 ;
        RECT 96.64 57.84 96.84 58.04 ;
        RECT 96.64 53.76 96.84 53.96 ;
        RECT 96.64 49.68 96.84 49.88 ;
        RECT 96.64 45.6 96.84 45.8 ;
        RECT 96.64 41.52 96.84 41.72 ;
        RECT 96.64 37.44 96.84 37.64 ;
        RECT 96.64 33.36 96.84 33.56 ;
        RECT 96.64 29.28 96.84 29.48 ;
        RECT 96.64 25.2 96.84 25.4 ;
        RECT 96.64 21.12 96.84 21.32 ;
        RECT 96.64 17.04 96.84 17.24 ;
        RECT 96.64 12.96 96.84 13.16 ;
        RECT 97.04 57.84 97.24 58.04 ;
        RECT 97.04 53.76 97.24 53.96 ;
        RECT 97.04 49.68 97.24 49.88 ;
        RECT 97.04 45.6 97.24 45.8 ;
        RECT 97.04 41.52 97.24 41.72 ;
        RECT 97.04 37.44 97.24 37.64 ;
        RECT 97.04 33.36 97.24 33.56 ;
        RECT 97.04 29.28 97.24 29.48 ;
        RECT 97.04 25.2 97.24 25.4 ;
        RECT 97.04 21.12 97.24 21.32 ;
        RECT 97.04 17.04 97.24 17.24 ;
        RECT 97.04 12.96 97.24 13.16 ;
        RECT 102.16 57.84 102.36 58.04 ;
        RECT 102.16 53.76 102.36 53.96 ;
        RECT 102.16 49.68 102.36 49.88 ;
        RECT 102.16 45.6 102.36 45.8 ;
        RECT 102.16 41.52 102.36 41.72 ;
        RECT 102.16 37.44 102.36 37.64 ;
        RECT 102.16 33.36 102.36 33.56 ;
        RECT 102.16 29.28 102.36 29.48 ;
        RECT 102.16 25.2 102.36 25.4 ;
        RECT 102.16 21.12 102.36 21.32 ;
        RECT 102.16 17.04 102.36 17.24 ;
        RECT 102.16 12.96 102.36 13.16 ;
        RECT 102.56 57.84 102.76 58.04 ;
        RECT 102.56 53.76 102.76 53.96 ;
        RECT 102.56 49.68 102.76 49.88 ;
        RECT 102.56 45.6 102.76 45.8 ;
        RECT 102.56 41.52 102.76 41.72 ;
        RECT 102.56 37.44 102.76 37.64 ;
        RECT 102.56 33.36 102.76 33.56 ;
        RECT 102.56 29.28 102.76 29.48 ;
        RECT 102.56 25.2 102.76 25.4 ;
        RECT 102.56 21.12 102.76 21.32 ;
        RECT 102.56 17.04 102.76 17.24 ;
        RECT 102.56 12.96 102.76 13.16 ;
        RECT 107.68 57.84 107.88 58.04 ;
        RECT 107.68 53.76 107.88 53.96 ;
        RECT 107.68 49.68 107.88 49.88 ;
        RECT 107.68 45.6 107.88 45.8 ;
        RECT 107.68 41.52 107.88 41.72 ;
        RECT 107.68 37.44 107.88 37.64 ;
        RECT 107.68 33.36 107.88 33.56 ;
        RECT 107.68 29.28 107.88 29.48 ;
        RECT 107.68 25.2 107.88 25.4 ;
        RECT 107.68 21.12 107.88 21.32 ;
        RECT 107.68 17.04 107.88 17.24 ;
        RECT 107.68 12.96 107.88 13.16 ;
        RECT 108.08 57.84 108.28 58.04 ;
        RECT 108.08 53.76 108.28 53.96 ;
        RECT 108.08 49.68 108.28 49.88 ;
        RECT 108.08 45.6 108.28 45.8 ;
        RECT 108.08 41.52 108.28 41.72 ;
        RECT 108.08 37.44 108.28 37.64 ;
        RECT 108.08 33.36 108.28 33.56 ;
        RECT 108.08 29.28 108.28 29.48 ;
        RECT 108.08 25.2 108.28 25.4 ;
        RECT 108.08 21.12 108.28 21.32 ;
        RECT 108.08 17.04 108.28 17.24 ;
        RECT 108.08 12.96 108.28 13.16 ;
        RECT 113.2 57.84 113.4 58.04 ;
        RECT 113.2 53.76 113.4 53.96 ;
        RECT 113.2 49.68 113.4 49.88 ;
        RECT 113.2 45.6 113.4 45.8 ;
        RECT 113.2 41.52 113.4 41.72 ;
        RECT 113.2 37.44 113.4 37.64 ;
        RECT 113.2 33.36 113.4 33.56 ;
        RECT 113.2 29.28 113.4 29.48 ;
        RECT 113.2 25.2 113.4 25.4 ;
        RECT 113.2 21.12 113.4 21.32 ;
        RECT 113.2 17.04 113.4 17.24 ;
        RECT 113.2 12.96 113.4 13.16 ;
        RECT 113.6 57.84 113.8 58.04 ;
        RECT 113.6 53.76 113.8 53.96 ;
        RECT 113.6 49.68 113.8 49.88 ;
        RECT 113.6 45.6 113.8 45.8 ;
        RECT 113.6 41.52 113.8 41.72 ;
        RECT 113.6 37.44 113.8 37.64 ;
        RECT 113.6 33.36 113.8 33.56 ;
        RECT 113.6 29.28 113.8 29.48 ;
        RECT 113.6 25.2 113.8 25.4 ;
        RECT 113.6 21.12 113.8 21.32 ;
        RECT 113.6 17.04 113.8 17.24 ;
        RECT 113.6 12.96 113.8 13.16 ;
        RECT 118.72 57.84 118.92 58.04 ;
        RECT 118.72 53.76 118.92 53.96 ;
        RECT 118.72 49.68 118.92 49.88 ;
        RECT 118.72 45.6 118.92 45.8 ;
        RECT 118.72 41.52 118.92 41.72 ;
        RECT 118.72 37.44 118.92 37.64 ;
        RECT 118.72 33.36 118.92 33.56 ;
        RECT 118.72 29.28 118.92 29.48 ;
        RECT 118.72 25.2 118.92 25.4 ;
        RECT 118.72 21.12 118.92 21.32 ;
        RECT 118.72 17.04 118.92 17.24 ;
        RECT 118.72 12.96 118.92 13.16 ;
        RECT 119.12 57.84 119.32 58.04 ;
        RECT 119.12 53.76 119.32 53.96 ;
        RECT 119.12 49.68 119.32 49.88 ;
        RECT 119.12 45.6 119.32 45.8 ;
        RECT 119.12 41.52 119.32 41.72 ;
        RECT 119.12 37.44 119.32 37.64 ;
        RECT 119.12 33.36 119.32 33.56 ;
        RECT 119.12 29.28 119.32 29.48 ;
        RECT 119.12 25.2 119.32 25.4 ;
        RECT 119.12 21.12 119.32 21.32 ;
        RECT 119.12 17.04 119.32 17.24 ;
        RECT 119.12 12.96 119.32 13.16 ;
        RECT 124.24 57.84 124.44 58.04 ;
        RECT 124.24 53.76 124.44 53.96 ;
        RECT 124.24 49.68 124.44 49.88 ;
        RECT 124.24 45.6 124.44 45.8 ;
        RECT 124.24 41.52 124.44 41.72 ;
        RECT 124.24 37.44 124.44 37.64 ;
        RECT 124.24 33.36 124.44 33.56 ;
        RECT 124.24 29.28 124.44 29.48 ;
        RECT 124.24 25.2 124.44 25.4 ;
        RECT 124.24 21.12 124.44 21.32 ;
        RECT 124.24 17.04 124.44 17.24 ;
        RECT 124.24 12.96 124.44 13.16 ;
        RECT 124.64 57.84 124.84 58.04 ;
        RECT 124.64 53.76 124.84 53.96 ;
        RECT 124.64 49.68 124.84 49.88 ;
        RECT 124.64 45.6 124.84 45.8 ;
        RECT 124.64 41.52 124.84 41.72 ;
        RECT 124.64 37.44 124.84 37.64 ;
        RECT 124.64 33.36 124.84 33.56 ;
        RECT 124.64 29.28 124.84 29.48 ;
        RECT 124.64 25.2 124.84 25.4 ;
        RECT 124.64 21.12 124.84 21.32 ;
        RECT 124.64 17.04 124.84 17.24 ;
        RECT 124.64 12.96 124.84 13.16 ;
        RECT 129.76 57.84 129.96 58.04 ;
        RECT 129.76 53.76 129.96 53.96 ;
        RECT 129.76 49.68 129.96 49.88 ;
        RECT 129.76 45.6 129.96 45.8 ;
        RECT 129.76 41.52 129.96 41.72 ;
        RECT 129.76 37.44 129.96 37.64 ;
        RECT 129.76 33.36 129.96 33.56 ;
        RECT 129.76 29.28 129.96 29.48 ;
        RECT 129.76 25.2 129.96 25.4 ;
        RECT 129.76 21.12 129.96 21.32 ;
        RECT 129.76 17.04 129.96 17.24 ;
        RECT 129.76 12.96 129.96 13.16 ;
        RECT 130.16 57.84 130.36 58.04 ;
        RECT 130.16 53.76 130.36 53.96 ;
        RECT 130.16 49.68 130.36 49.88 ;
        RECT 130.16 45.6 130.36 45.8 ;
        RECT 130.16 41.52 130.36 41.72 ;
        RECT 130.16 37.44 130.36 37.64 ;
        RECT 130.16 33.36 130.36 33.56 ;
        RECT 130.16 29.28 130.36 29.48 ;
        RECT 130.16 25.2 130.36 25.4 ;
        RECT 130.16 21.12 130.36 21.32 ;
        RECT 130.16 17.04 130.36 17.24 ;
        RECT 130.16 12.96 130.36 13.16 ;
        RECT 135.28 57.84 135.48 58.04 ;
        RECT 135.28 53.76 135.48 53.96 ;
        RECT 135.28 49.68 135.48 49.88 ;
        RECT 135.28 45.6 135.48 45.8 ;
        RECT 135.28 41.52 135.48 41.72 ;
        RECT 135.28 37.44 135.48 37.64 ;
        RECT 135.28 33.36 135.48 33.56 ;
        RECT 135.28 29.28 135.48 29.48 ;
        RECT 135.28 25.2 135.48 25.4 ;
        RECT 135.28 21.12 135.48 21.32 ;
        RECT 135.28 17.04 135.48 17.24 ;
        RECT 135.28 12.96 135.48 13.16 ;
        RECT 135.68 57.84 135.88 58.04 ;
        RECT 135.68 53.76 135.88 53.96 ;
        RECT 135.68 49.68 135.88 49.88 ;
        RECT 135.68 45.6 135.88 45.8 ;
        RECT 135.68 41.52 135.88 41.72 ;
        RECT 135.68 37.44 135.88 37.64 ;
        RECT 135.68 33.36 135.88 33.56 ;
        RECT 135.68 29.28 135.88 29.48 ;
        RECT 135.68 25.2 135.88 25.4 ;
        RECT 135.68 21.12 135.88 21.32 ;
        RECT 135.68 17.04 135.88 17.24 ;
        RECT 135.68 12.96 135.88 13.16 ;
        RECT 140.8 57.84 141 58.04 ;
        RECT 140.8 53.76 141 53.96 ;
        RECT 140.8 49.68 141 49.88 ;
        RECT 140.8 45.6 141 45.8 ;
        RECT 140.8 41.52 141 41.72 ;
        RECT 140.8 37.44 141 37.64 ;
        RECT 140.8 33.36 141 33.56 ;
        RECT 140.8 29.28 141 29.48 ;
        RECT 140.8 25.2 141 25.4 ;
        RECT 140.8 21.12 141 21.32 ;
        RECT 140.8 17.04 141 17.24 ;
        RECT 140.8 12.96 141 13.16 ;
        RECT 141.2 57.84 141.4 58.04 ;
        RECT 141.2 53.76 141.4 53.96 ;
        RECT 141.2 49.68 141.4 49.88 ;
        RECT 141.2 45.6 141.4 45.8 ;
        RECT 141.2 41.52 141.4 41.72 ;
        RECT 141.2 37.44 141.4 37.64 ;
        RECT 141.2 33.36 141.4 33.56 ;
        RECT 141.2 29.28 141.4 29.48 ;
        RECT 141.2 25.2 141.4 25.4 ;
        RECT 141.2 21.12 141.4 21.32 ;
        RECT 141.2 17.04 141.4 17.24 ;
        RECT 141.2 12.96 141.4 13.16 ;
        RECT 146.32 57.84 146.52 58.04 ;
        RECT 146.32 53.76 146.52 53.96 ;
        RECT 146.32 49.68 146.52 49.88 ;
        RECT 146.32 45.6 146.52 45.8 ;
        RECT 146.32 41.52 146.52 41.72 ;
        RECT 146.32 37.44 146.52 37.64 ;
        RECT 146.32 33.36 146.52 33.56 ;
        RECT 146.32 29.28 146.52 29.48 ;
        RECT 146.32 25.2 146.52 25.4 ;
        RECT 146.32 21.12 146.52 21.32 ;
        RECT 146.32 17.04 146.52 17.24 ;
        RECT 146.32 12.96 146.52 13.16 ;
        RECT 146.72 57.84 146.92 58.04 ;
        RECT 146.72 53.76 146.92 53.96 ;
        RECT 146.72 49.68 146.92 49.88 ;
        RECT 146.72 45.6 146.92 45.8 ;
        RECT 146.72 41.52 146.92 41.72 ;
        RECT 146.72 37.44 146.92 37.64 ;
        RECT 146.72 33.36 146.92 33.56 ;
        RECT 146.72 29.28 146.92 29.48 ;
        RECT 146.72 25.2 146.92 25.4 ;
        RECT 146.72 21.12 146.92 21.32 ;
        RECT 146.72 17.04 146.92 17.24 ;
        RECT 146.72 12.96 146.92 13.16 ;
        RECT 151.84 57.84 152.04 58.04 ;
        RECT 151.84 53.76 152.04 53.96 ;
        RECT 151.84 49.68 152.04 49.88 ;
        RECT 151.84 45.6 152.04 45.8 ;
        RECT 151.84 41.52 152.04 41.72 ;
        RECT 151.84 37.44 152.04 37.64 ;
        RECT 151.84 33.36 152.04 33.56 ;
        RECT 151.84 29.28 152.04 29.48 ;
        RECT 151.84 25.2 152.04 25.4 ;
        RECT 151.84 21.12 152.04 21.32 ;
        RECT 151.84 17.04 152.04 17.24 ;
        RECT 151.84 12.96 152.04 13.16 ;
        RECT 152.24 57.84 152.44 58.04 ;
        RECT 152.24 53.76 152.44 53.96 ;
        RECT 152.24 49.68 152.44 49.88 ;
        RECT 152.24 45.6 152.44 45.8 ;
        RECT 152.24 41.52 152.44 41.72 ;
        RECT 152.24 37.44 152.44 37.64 ;
        RECT 152.24 33.36 152.44 33.56 ;
        RECT 152.24 29.28 152.44 29.48 ;
        RECT 152.24 25.2 152.44 25.4 ;
        RECT 152.24 21.12 152.44 21.32 ;
        RECT 152.24 17.04 152.44 17.24 ;
        RECT 152.24 12.96 152.44 13.16 ;
        RECT 157.36 57.84 157.56 58.04 ;
        RECT 157.36 53.76 157.56 53.96 ;
        RECT 157.36 49.68 157.56 49.88 ;
        RECT 157.36 45.6 157.56 45.8 ;
        RECT 157.36 41.52 157.56 41.72 ;
        RECT 157.36 37.44 157.56 37.64 ;
        RECT 157.36 33.36 157.56 33.56 ;
        RECT 157.36 29.28 157.56 29.48 ;
        RECT 157.36 25.2 157.56 25.4 ;
        RECT 157.36 21.12 157.56 21.32 ;
        RECT 157.36 17.04 157.56 17.24 ;
        RECT 157.36 12.96 157.56 13.16 ;
        RECT 157.76 57.84 157.96 58.04 ;
        RECT 157.76 53.76 157.96 53.96 ;
        RECT 157.76 49.68 157.96 49.88 ;
        RECT 157.76 45.6 157.96 45.8 ;
        RECT 157.76 41.52 157.96 41.72 ;
        RECT 157.76 37.44 157.96 37.64 ;
        RECT 157.76 33.36 157.96 33.56 ;
        RECT 157.76 29.28 157.96 29.48 ;
        RECT 157.76 25.2 157.96 25.4 ;
        RECT 157.76 21.12 157.96 21.32 ;
        RECT 157.76 17.04 157.96 17.24 ;
        RECT 157.76 12.96 157.96 13.16 ;
        RECT 162.88 57.84 163.08 58.04 ;
        RECT 162.88 53.76 163.08 53.96 ;
        RECT 162.88 49.68 163.08 49.88 ;
        RECT 162.88 45.6 163.08 45.8 ;
        RECT 162.88 41.52 163.08 41.72 ;
        RECT 162.88 37.44 163.08 37.64 ;
        RECT 162.88 33.36 163.08 33.56 ;
        RECT 162.88 29.28 163.08 29.48 ;
        RECT 162.88 25.2 163.08 25.4 ;
        RECT 162.88 21.12 163.08 21.32 ;
        RECT 162.88 17.04 163.08 17.24 ;
        RECT 162.88 12.96 163.08 13.16 ;
        RECT 163.28 57.84 163.48 58.04 ;
        RECT 163.28 53.76 163.48 53.96 ;
        RECT 163.28 49.68 163.48 49.88 ;
        RECT 163.28 45.6 163.48 45.8 ;
        RECT 163.28 41.52 163.48 41.72 ;
        RECT 163.28 37.44 163.48 37.64 ;
        RECT 163.28 33.36 163.48 33.56 ;
        RECT 163.28 29.28 163.48 29.48 ;
        RECT 163.28 25.2 163.48 25.4 ;
        RECT 163.28 21.12 163.48 21.32 ;
        RECT 163.28 17.04 163.48 17.24 ;
        RECT 163.28 12.96 163.48 13.16 ;
        RECT 168.4 57.84 168.6 58.04 ;
        RECT 168.4 53.76 168.6 53.96 ;
        RECT 168.4 49.68 168.6 49.88 ;
        RECT 168.4 45.6 168.6 45.8 ;
        RECT 168.4 41.52 168.6 41.72 ;
        RECT 168.4 37.44 168.6 37.64 ;
        RECT 168.4 33.36 168.6 33.56 ;
        RECT 168.4 29.28 168.6 29.48 ;
        RECT 168.4 25.2 168.6 25.4 ;
        RECT 168.4 21.12 168.6 21.32 ;
        RECT 168.4 17.04 168.6 17.24 ;
        RECT 168.4 12.96 168.6 13.16 ;
        RECT 168.8 57.84 169 58.04 ;
        RECT 168.8 53.76 169 53.96 ;
        RECT 168.8 49.68 169 49.88 ;
        RECT 168.8 45.6 169 45.8 ;
        RECT 168.8 41.52 169 41.72 ;
        RECT 168.8 37.44 169 37.64 ;
        RECT 168.8 33.36 169 33.56 ;
        RECT 168.8 29.28 169 29.48 ;
        RECT 168.8 25.2 169 25.4 ;
        RECT 168.8 21.12 169 21.32 ;
        RECT 168.8 17.04 169 17.24 ;
        RECT 168.8 12.96 169 13.16 ;
        RECT 173.92 57.84 174.12 58.04 ;
        RECT 173.92 53.76 174.12 53.96 ;
        RECT 173.92 49.68 174.12 49.88 ;
        RECT 173.92 45.6 174.12 45.8 ;
        RECT 173.92 41.52 174.12 41.72 ;
        RECT 173.92 37.44 174.12 37.64 ;
        RECT 173.92 33.36 174.12 33.56 ;
        RECT 173.92 29.28 174.12 29.48 ;
        RECT 173.92 25.2 174.12 25.4 ;
        RECT 173.92 21.12 174.12 21.32 ;
        RECT 173.92 17.04 174.12 17.24 ;
        RECT 173.92 12.96 174.12 13.16 ;
        RECT 174.32 57.84 174.52 58.04 ;
        RECT 174.32 53.76 174.52 53.96 ;
        RECT 174.32 49.68 174.52 49.88 ;
        RECT 174.32 45.6 174.52 45.8 ;
        RECT 174.32 41.52 174.52 41.72 ;
        RECT 174.32 37.44 174.52 37.64 ;
        RECT 174.32 33.36 174.52 33.56 ;
        RECT 174.32 29.28 174.52 29.48 ;
        RECT 174.32 25.2 174.52 25.4 ;
        RECT 174.32 21.12 174.52 21.32 ;
        RECT 174.32 17.04 174.52 17.24 ;
        RECT 174.32 12.96 174.52 13.16 ;
        RECT 179.44 57.84 179.64 58.04 ;
        RECT 179.44 53.76 179.64 53.96 ;
        RECT 179.44 49.68 179.64 49.88 ;
        RECT 179.44 45.6 179.64 45.8 ;
        RECT 179.44 41.52 179.64 41.72 ;
        RECT 179.44 37.44 179.64 37.64 ;
        RECT 179.44 33.36 179.64 33.56 ;
        RECT 179.44 29.28 179.64 29.48 ;
        RECT 179.44 25.2 179.64 25.4 ;
        RECT 179.44 21.12 179.64 21.32 ;
        RECT 179.44 17.04 179.64 17.24 ;
        RECT 179.44 12.96 179.64 13.16 ;
        RECT 179.84 57.84 180.04 58.04 ;
        RECT 179.84 53.76 180.04 53.96 ;
        RECT 179.84 49.68 180.04 49.88 ;
        RECT 179.84 45.6 180.04 45.8 ;
        RECT 179.84 41.52 180.04 41.72 ;
        RECT 179.84 37.44 180.04 37.64 ;
        RECT 179.84 33.36 180.04 33.56 ;
        RECT 179.84 29.28 180.04 29.48 ;
        RECT 179.84 25.2 180.04 25.4 ;
        RECT 179.84 21.12 180.04 21.32 ;
        RECT 179.84 17.04 180.04 17.24 ;
        RECT 179.84 12.96 180.04 13.16 ;
        RECT 184.96 57.84 185.16 58.04 ;
        RECT 184.96 53.76 185.16 53.96 ;
        RECT 184.96 49.68 185.16 49.88 ;
        RECT 184.96 45.6 185.16 45.8 ;
        RECT 184.96 41.52 185.16 41.72 ;
        RECT 184.96 37.44 185.16 37.64 ;
        RECT 184.96 33.36 185.16 33.56 ;
        RECT 184.96 29.28 185.16 29.48 ;
        RECT 184.96 25.2 185.16 25.4 ;
        RECT 184.96 21.12 185.16 21.32 ;
        RECT 184.96 17.04 185.16 17.24 ;
        RECT 184.96 12.96 185.16 13.16 ;
        RECT 185.36 57.84 185.56 58.04 ;
        RECT 185.36 53.76 185.56 53.96 ;
        RECT 185.36 49.68 185.56 49.88 ;
        RECT 185.36 45.6 185.56 45.8 ;
        RECT 185.36 41.52 185.56 41.72 ;
        RECT 185.36 37.44 185.56 37.64 ;
        RECT 185.36 33.36 185.56 33.56 ;
        RECT 185.36 29.28 185.56 29.48 ;
        RECT 185.36 25.2 185.56 25.4 ;
        RECT 185.36 21.12 185.56 21.32 ;
        RECT 185.36 17.04 185.56 17.24 ;
        RECT 185.36 12.96 185.56 13.16 ;
      LAYER via ;
        RECT 11.995 58.885 12.145 59.035 ;
        RECT 11.995 53.445 12.145 53.595 ;
        RECT 11.995 48.005 12.145 48.155 ;
        RECT 11.995 42.565 12.145 42.715 ;
        RECT 11.995 37.125 12.145 37.275 ;
        RECT 11.995 31.685 12.145 31.835 ;
        RECT 11.995 26.245 12.145 26.395 ;
        RECT 11.995 20.805 12.145 20.955 ;
        RECT 11.995 15.365 12.145 15.515 ;
        RECT 11.995 10.035 12.145 10.185 ;
        RECT 14.755 58.885 14.905 59.035 ;
        RECT 14.755 53.445 14.905 53.595 ;
        RECT 14.755 48.005 14.905 48.155 ;
        RECT 14.755 42.565 14.905 42.715 ;
        RECT 14.755 37.125 14.905 37.275 ;
        RECT 14.755 31.685 14.905 31.835 ;
        RECT 14.755 26.245 14.905 26.395 ;
        RECT 14.755 20.805 14.905 20.955 ;
        RECT 14.755 15.365 14.905 15.515 ;
        RECT 14.755 10.035 14.905 10.185 ;
        RECT 17.515 58.885 17.665 59.035 ;
        RECT 17.515 53.445 17.665 53.595 ;
        RECT 17.515 48.005 17.665 48.155 ;
        RECT 17.515 42.565 17.665 42.715 ;
        RECT 17.515 37.125 17.665 37.275 ;
        RECT 17.515 31.685 17.665 31.835 ;
        RECT 17.515 26.245 17.665 26.395 ;
        RECT 17.515 20.805 17.665 20.955 ;
        RECT 17.515 15.365 17.665 15.515 ;
        RECT 17.515 10.035 17.665 10.185 ;
        RECT 20.275 58.885 20.425 59.035 ;
        RECT 20.275 53.445 20.425 53.595 ;
        RECT 20.275 48.005 20.425 48.155 ;
        RECT 20.275 42.565 20.425 42.715 ;
        RECT 20.275 37.125 20.425 37.275 ;
        RECT 20.275 31.685 20.425 31.835 ;
        RECT 20.275 26.245 20.425 26.395 ;
        RECT 20.275 20.805 20.425 20.955 ;
        RECT 20.275 15.365 20.425 15.515 ;
        RECT 20.275 10.035 20.425 10.185 ;
        RECT 23.035 58.885 23.185 59.035 ;
        RECT 23.035 53.445 23.185 53.595 ;
        RECT 23.035 48.005 23.185 48.155 ;
        RECT 23.035 42.565 23.185 42.715 ;
        RECT 23.035 37.125 23.185 37.275 ;
        RECT 23.035 31.685 23.185 31.835 ;
        RECT 23.035 26.245 23.185 26.395 ;
        RECT 23.035 20.805 23.185 20.955 ;
        RECT 23.035 15.365 23.185 15.515 ;
        RECT 23.035 10.035 23.185 10.185 ;
        RECT 25.795 58.885 25.945 59.035 ;
        RECT 25.795 53.445 25.945 53.595 ;
        RECT 25.795 48.005 25.945 48.155 ;
        RECT 25.795 42.565 25.945 42.715 ;
        RECT 25.795 37.125 25.945 37.275 ;
        RECT 25.795 31.685 25.945 31.835 ;
        RECT 25.795 26.245 25.945 26.395 ;
        RECT 25.795 20.805 25.945 20.955 ;
        RECT 25.795 15.365 25.945 15.515 ;
        RECT 25.795 10.035 25.945 10.185 ;
        RECT 28.555 58.885 28.705 59.035 ;
        RECT 28.555 53.445 28.705 53.595 ;
        RECT 28.555 48.005 28.705 48.155 ;
        RECT 28.555 42.565 28.705 42.715 ;
        RECT 28.555 37.125 28.705 37.275 ;
        RECT 28.555 31.685 28.705 31.835 ;
        RECT 28.555 26.245 28.705 26.395 ;
        RECT 28.555 20.805 28.705 20.955 ;
        RECT 28.555 15.365 28.705 15.515 ;
        RECT 28.555 10.035 28.705 10.185 ;
        RECT 31.315 58.885 31.465 59.035 ;
        RECT 31.315 53.445 31.465 53.595 ;
        RECT 31.315 48.005 31.465 48.155 ;
        RECT 31.315 42.565 31.465 42.715 ;
        RECT 31.315 37.125 31.465 37.275 ;
        RECT 31.315 31.685 31.465 31.835 ;
        RECT 31.315 26.245 31.465 26.395 ;
        RECT 31.315 20.805 31.465 20.955 ;
        RECT 31.315 15.365 31.465 15.515 ;
        RECT 31.315 10.035 31.465 10.185 ;
        RECT 34.075 58.885 34.225 59.035 ;
        RECT 34.075 53.445 34.225 53.595 ;
        RECT 34.075 48.005 34.225 48.155 ;
        RECT 34.075 42.565 34.225 42.715 ;
        RECT 34.075 37.125 34.225 37.275 ;
        RECT 34.075 31.685 34.225 31.835 ;
        RECT 34.075 26.245 34.225 26.395 ;
        RECT 34.075 20.805 34.225 20.955 ;
        RECT 34.075 15.365 34.225 15.515 ;
        RECT 34.075 10.035 34.225 10.185 ;
        RECT 36.835 58.885 36.985 59.035 ;
        RECT 36.835 53.445 36.985 53.595 ;
        RECT 36.835 48.005 36.985 48.155 ;
        RECT 36.835 42.565 36.985 42.715 ;
        RECT 36.835 37.125 36.985 37.275 ;
        RECT 36.835 31.685 36.985 31.835 ;
        RECT 36.835 26.245 36.985 26.395 ;
        RECT 36.835 20.805 36.985 20.955 ;
        RECT 36.835 15.365 36.985 15.515 ;
        RECT 36.835 10.035 36.985 10.185 ;
        RECT 39.595 58.885 39.745 59.035 ;
        RECT 39.595 53.445 39.745 53.595 ;
        RECT 39.595 48.005 39.745 48.155 ;
        RECT 39.595 42.565 39.745 42.715 ;
        RECT 39.595 37.125 39.745 37.275 ;
        RECT 39.595 31.685 39.745 31.835 ;
        RECT 39.595 26.245 39.745 26.395 ;
        RECT 39.595 20.805 39.745 20.955 ;
        RECT 39.595 15.365 39.745 15.515 ;
        RECT 39.595 10.035 39.745 10.185 ;
        RECT 42.355 58.885 42.505 59.035 ;
        RECT 42.355 53.445 42.505 53.595 ;
        RECT 42.355 48.005 42.505 48.155 ;
        RECT 42.355 42.565 42.505 42.715 ;
        RECT 42.355 37.125 42.505 37.275 ;
        RECT 42.355 31.685 42.505 31.835 ;
        RECT 42.355 26.245 42.505 26.395 ;
        RECT 42.355 20.805 42.505 20.955 ;
        RECT 42.355 15.365 42.505 15.515 ;
        RECT 42.355 10.035 42.505 10.185 ;
        RECT 45.115 58.885 45.265 59.035 ;
        RECT 45.115 53.445 45.265 53.595 ;
        RECT 45.115 48.005 45.265 48.155 ;
        RECT 45.115 42.565 45.265 42.715 ;
        RECT 45.115 37.125 45.265 37.275 ;
        RECT 45.115 31.685 45.265 31.835 ;
        RECT 45.115 26.245 45.265 26.395 ;
        RECT 45.115 20.805 45.265 20.955 ;
        RECT 45.115 15.365 45.265 15.515 ;
        RECT 45.115 10.035 45.265 10.185 ;
        RECT 47.875 58.885 48.025 59.035 ;
        RECT 47.875 53.445 48.025 53.595 ;
        RECT 47.875 48.005 48.025 48.155 ;
        RECT 47.875 42.565 48.025 42.715 ;
        RECT 47.875 37.125 48.025 37.275 ;
        RECT 47.875 31.685 48.025 31.835 ;
        RECT 47.875 26.245 48.025 26.395 ;
        RECT 47.875 20.805 48.025 20.955 ;
        RECT 47.875 15.365 48.025 15.515 ;
        RECT 47.875 10.035 48.025 10.185 ;
        RECT 50.635 58.885 50.785 59.035 ;
        RECT 50.635 53.445 50.785 53.595 ;
        RECT 50.635 48.005 50.785 48.155 ;
        RECT 50.635 42.565 50.785 42.715 ;
        RECT 50.635 37.125 50.785 37.275 ;
        RECT 50.635 31.685 50.785 31.835 ;
        RECT 50.635 26.245 50.785 26.395 ;
        RECT 50.635 20.805 50.785 20.955 ;
        RECT 50.635 15.365 50.785 15.515 ;
        RECT 50.635 10.035 50.785 10.185 ;
        RECT 53.395 58.885 53.545 59.035 ;
        RECT 53.395 53.445 53.545 53.595 ;
        RECT 53.395 48.005 53.545 48.155 ;
        RECT 53.395 42.565 53.545 42.715 ;
        RECT 53.395 37.125 53.545 37.275 ;
        RECT 53.395 31.685 53.545 31.835 ;
        RECT 53.395 26.245 53.545 26.395 ;
        RECT 53.395 20.805 53.545 20.955 ;
        RECT 53.395 15.365 53.545 15.515 ;
        RECT 53.395 10.035 53.545 10.185 ;
        RECT 56.155 58.885 56.305 59.035 ;
        RECT 56.155 53.445 56.305 53.595 ;
        RECT 56.155 48.005 56.305 48.155 ;
        RECT 56.155 42.565 56.305 42.715 ;
        RECT 56.155 37.125 56.305 37.275 ;
        RECT 56.155 31.685 56.305 31.835 ;
        RECT 56.155 26.245 56.305 26.395 ;
        RECT 56.155 20.805 56.305 20.955 ;
        RECT 56.155 15.365 56.305 15.515 ;
        RECT 56.155 10.035 56.305 10.185 ;
        RECT 58.915 58.885 59.065 59.035 ;
        RECT 58.915 53.445 59.065 53.595 ;
        RECT 58.915 48.005 59.065 48.155 ;
        RECT 58.915 42.565 59.065 42.715 ;
        RECT 58.915 37.125 59.065 37.275 ;
        RECT 58.915 31.685 59.065 31.835 ;
        RECT 58.915 26.245 59.065 26.395 ;
        RECT 58.915 20.805 59.065 20.955 ;
        RECT 58.915 15.365 59.065 15.515 ;
        RECT 58.915 10.035 59.065 10.185 ;
        RECT 61.675 58.885 61.825 59.035 ;
        RECT 61.675 53.445 61.825 53.595 ;
        RECT 61.675 48.005 61.825 48.155 ;
        RECT 61.675 42.565 61.825 42.715 ;
        RECT 61.675 37.125 61.825 37.275 ;
        RECT 61.675 31.685 61.825 31.835 ;
        RECT 61.675 26.245 61.825 26.395 ;
        RECT 61.675 20.805 61.825 20.955 ;
        RECT 61.675 15.365 61.825 15.515 ;
        RECT 61.675 10.035 61.825 10.185 ;
        RECT 64.435 58.885 64.585 59.035 ;
        RECT 64.435 53.445 64.585 53.595 ;
        RECT 64.435 48.005 64.585 48.155 ;
        RECT 64.435 42.565 64.585 42.715 ;
        RECT 64.435 37.125 64.585 37.275 ;
        RECT 64.435 31.685 64.585 31.835 ;
        RECT 64.435 26.245 64.585 26.395 ;
        RECT 64.435 20.805 64.585 20.955 ;
        RECT 64.435 15.365 64.585 15.515 ;
        RECT 64.435 10.035 64.585 10.185 ;
        RECT 67.195 58.885 67.345 59.035 ;
        RECT 67.195 53.445 67.345 53.595 ;
        RECT 67.195 48.005 67.345 48.155 ;
        RECT 67.195 42.565 67.345 42.715 ;
        RECT 67.195 37.125 67.345 37.275 ;
        RECT 67.195 31.685 67.345 31.835 ;
        RECT 67.195 26.245 67.345 26.395 ;
        RECT 67.195 20.805 67.345 20.955 ;
        RECT 67.195 15.365 67.345 15.515 ;
        RECT 67.195 10.035 67.345 10.185 ;
        RECT 69.955 58.885 70.105 59.035 ;
        RECT 69.955 53.445 70.105 53.595 ;
        RECT 69.955 48.005 70.105 48.155 ;
        RECT 69.955 42.565 70.105 42.715 ;
        RECT 69.955 37.125 70.105 37.275 ;
        RECT 69.955 31.685 70.105 31.835 ;
        RECT 69.955 26.245 70.105 26.395 ;
        RECT 69.955 20.805 70.105 20.955 ;
        RECT 69.955 15.365 70.105 15.515 ;
        RECT 69.955 10.035 70.105 10.185 ;
        RECT 72.715 58.885 72.865 59.035 ;
        RECT 72.715 53.445 72.865 53.595 ;
        RECT 72.715 48.005 72.865 48.155 ;
        RECT 72.715 42.565 72.865 42.715 ;
        RECT 72.715 37.125 72.865 37.275 ;
        RECT 72.715 31.685 72.865 31.835 ;
        RECT 72.715 26.245 72.865 26.395 ;
        RECT 72.715 20.805 72.865 20.955 ;
        RECT 72.715 15.365 72.865 15.515 ;
        RECT 72.715 10.035 72.865 10.185 ;
        RECT 75.475 58.885 75.625 59.035 ;
        RECT 75.475 53.445 75.625 53.595 ;
        RECT 75.475 48.005 75.625 48.155 ;
        RECT 75.475 42.565 75.625 42.715 ;
        RECT 75.475 37.125 75.625 37.275 ;
        RECT 75.475 31.685 75.625 31.835 ;
        RECT 75.475 26.245 75.625 26.395 ;
        RECT 75.475 20.805 75.625 20.955 ;
        RECT 75.475 15.365 75.625 15.515 ;
        RECT 75.475 10.035 75.625 10.185 ;
        RECT 78.235 58.885 78.385 59.035 ;
        RECT 78.235 53.445 78.385 53.595 ;
        RECT 78.235 48.005 78.385 48.155 ;
        RECT 78.235 42.565 78.385 42.715 ;
        RECT 78.235 37.125 78.385 37.275 ;
        RECT 78.235 31.685 78.385 31.835 ;
        RECT 78.235 26.245 78.385 26.395 ;
        RECT 78.235 20.805 78.385 20.955 ;
        RECT 78.235 15.365 78.385 15.515 ;
        RECT 78.235 10.035 78.385 10.185 ;
        RECT 80.995 58.885 81.145 59.035 ;
        RECT 80.995 53.445 81.145 53.595 ;
        RECT 80.995 48.005 81.145 48.155 ;
        RECT 80.995 42.565 81.145 42.715 ;
        RECT 80.995 37.125 81.145 37.275 ;
        RECT 80.995 31.685 81.145 31.835 ;
        RECT 80.995 26.245 81.145 26.395 ;
        RECT 80.995 20.805 81.145 20.955 ;
        RECT 80.995 15.365 81.145 15.515 ;
        RECT 80.995 10.035 81.145 10.185 ;
        RECT 83.755 58.885 83.905 59.035 ;
        RECT 83.755 53.445 83.905 53.595 ;
        RECT 83.755 48.005 83.905 48.155 ;
        RECT 83.755 42.565 83.905 42.715 ;
        RECT 83.755 37.125 83.905 37.275 ;
        RECT 83.755 31.685 83.905 31.835 ;
        RECT 83.755 26.245 83.905 26.395 ;
        RECT 83.755 20.805 83.905 20.955 ;
        RECT 83.755 15.365 83.905 15.515 ;
        RECT 83.755 10.035 83.905 10.185 ;
        RECT 86.515 58.885 86.665 59.035 ;
        RECT 86.515 53.445 86.665 53.595 ;
        RECT 86.515 48.005 86.665 48.155 ;
        RECT 86.515 42.565 86.665 42.715 ;
        RECT 86.515 37.125 86.665 37.275 ;
        RECT 86.515 31.685 86.665 31.835 ;
        RECT 86.515 26.245 86.665 26.395 ;
        RECT 86.515 20.805 86.665 20.955 ;
        RECT 86.515 15.365 86.665 15.515 ;
        RECT 86.515 10.035 86.665 10.185 ;
        RECT 89.275 58.885 89.425 59.035 ;
        RECT 89.275 53.445 89.425 53.595 ;
        RECT 89.275 48.005 89.425 48.155 ;
        RECT 89.275 42.565 89.425 42.715 ;
        RECT 89.275 37.125 89.425 37.275 ;
        RECT 89.275 31.685 89.425 31.835 ;
        RECT 89.275 26.245 89.425 26.395 ;
        RECT 89.275 20.805 89.425 20.955 ;
        RECT 89.275 15.365 89.425 15.515 ;
        RECT 89.275 10.035 89.425 10.185 ;
        RECT 92.035 58.885 92.185 59.035 ;
        RECT 92.035 53.445 92.185 53.595 ;
        RECT 92.035 48.005 92.185 48.155 ;
        RECT 92.035 42.565 92.185 42.715 ;
        RECT 92.035 37.125 92.185 37.275 ;
        RECT 92.035 31.685 92.185 31.835 ;
        RECT 92.035 26.245 92.185 26.395 ;
        RECT 92.035 20.805 92.185 20.955 ;
        RECT 92.035 15.365 92.185 15.515 ;
        RECT 92.035 10.035 92.185 10.185 ;
        RECT 94.795 58.885 94.945 59.035 ;
        RECT 94.795 53.445 94.945 53.595 ;
        RECT 94.795 48.005 94.945 48.155 ;
        RECT 94.795 42.565 94.945 42.715 ;
        RECT 94.795 37.125 94.945 37.275 ;
        RECT 94.795 31.685 94.945 31.835 ;
        RECT 94.795 26.245 94.945 26.395 ;
        RECT 94.795 20.805 94.945 20.955 ;
        RECT 94.795 15.365 94.945 15.515 ;
        RECT 94.795 10.035 94.945 10.185 ;
        RECT 97.555 58.885 97.705 59.035 ;
        RECT 97.555 53.445 97.705 53.595 ;
        RECT 97.555 48.005 97.705 48.155 ;
        RECT 97.555 42.565 97.705 42.715 ;
        RECT 97.555 37.125 97.705 37.275 ;
        RECT 97.555 31.685 97.705 31.835 ;
        RECT 97.555 26.245 97.705 26.395 ;
        RECT 97.555 20.805 97.705 20.955 ;
        RECT 97.555 15.365 97.705 15.515 ;
        RECT 97.555 10.035 97.705 10.185 ;
        RECT 100.315 58.885 100.465 59.035 ;
        RECT 100.315 53.445 100.465 53.595 ;
        RECT 100.315 48.005 100.465 48.155 ;
        RECT 100.315 42.565 100.465 42.715 ;
        RECT 100.315 37.125 100.465 37.275 ;
        RECT 100.315 31.685 100.465 31.835 ;
        RECT 100.315 26.245 100.465 26.395 ;
        RECT 100.315 20.805 100.465 20.955 ;
        RECT 100.315 15.365 100.465 15.515 ;
        RECT 100.315 10.035 100.465 10.185 ;
        RECT 103.075 58.885 103.225 59.035 ;
        RECT 103.075 53.445 103.225 53.595 ;
        RECT 103.075 48.005 103.225 48.155 ;
        RECT 103.075 42.565 103.225 42.715 ;
        RECT 103.075 37.125 103.225 37.275 ;
        RECT 103.075 31.685 103.225 31.835 ;
        RECT 103.075 26.245 103.225 26.395 ;
        RECT 103.075 20.805 103.225 20.955 ;
        RECT 103.075 15.365 103.225 15.515 ;
        RECT 103.075 10.035 103.225 10.185 ;
        RECT 105.835 58.885 105.985 59.035 ;
        RECT 105.835 53.445 105.985 53.595 ;
        RECT 105.835 48.005 105.985 48.155 ;
        RECT 105.835 42.565 105.985 42.715 ;
        RECT 105.835 37.125 105.985 37.275 ;
        RECT 105.835 31.685 105.985 31.835 ;
        RECT 105.835 26.245 105.985 26.395 ;
        RECT 105.835 20.805 105.985 20.955 ;
        RECT 105.835 15.365 105.985 15.515 ;
        RECT 105.835 10.035 105.985 10.185 ;
        RECT 108.595 58.885 108.745 59.035 ;
        RECT 108.595 53.445 108.745 53.595 ;
        RECT 108.595 48.005 108.745 48.155 ;
        RECT 108.595 42.565 108.745 42.715 ;
        RECT 108.595 37.125 108.745 37.275 ;
        RECT 108.595 31.685 108.745 31.835 ;
        RECT 108.595 26.245 108.745 26.395 ;
        RECT 108.595 20.805 108.745 20.955 ;
        RECT 108.595 15.365 108.745 15.515 ;
        RECT 108.595 10.035 108.745 10.185 ;
        RECT 111.355 58.885 111.505 59.035 ;
        RECT 111.355 53.445 111.505 53.595 ;
        RECT 111.355 48.005 111.505 48.155 ;
        RECT 111.355 42.565 111.505 42.715 ;
        RECT 111.355 37.125 111.505 37.275 ;
        RECT 111.355 31.685 111.505 31.835 ;
        RECT 111.355 26.245 111.505 26.395 ;
        RECT 111.355 20.805 111.505 20.955 ;
        RECT 111.355 15.365 111.505 15.515 ;
        RECT 111.355 10.035 111.505 10.185 ;
        RECT 114.115 58.885 114.265 59.035 ;
        RECT 114.115 53.445 114.265 53.595 ;
        RECT 114.115 48.005 114.265 48.155 ;
        RECT 114.115 42.565 114.265 42.715 ;
        RECT 114.115 37.125 114.265 37.275 ;
        RECT 114.115 31.685 114.265 31.835 ;
        RECT 114.115 26.245 114.265 26.395 ;
        RECT 114.115 20.805 114.265 20.955 ;
        RECT 114.115 15.365 114.265 15.515 ;
        RECT 114.115 10.035 114.265 10.185 ;
        RECT 116.875 58.885 117.025 59.035 ;
        RECT 116.875 53.445 117.025 53.595 ;
        RECT 116.875 48.005 117.025 48.155 ;
        RECT 116.875 42.565 117.025 42.715 ;
        RECT 116.875 37.125 117.025 37.275 ;
        RECT 116.875 31.685 117.025 31.835 ;
        RECT 116.875 26.245 117.025 26.395 ;
        RECT 116.875 20.805 117.025 20.955 ;
        RECT 116.875 15.365 117.025 15.515 ;
        RECT 116.875 10.035 117.025 10.185 ;
        RECT 119.635 58.885 119.785 59.035 ;
        RECT 119.635 53.445 119.785 53.595 ;
        RECT 119.635 48.005 119.785 48.155 ;
        RECT 119.635 42.565 119.785 42.715 ;
        RECT 119.635 37.125 119.785 37.275 ;
        RECT 119.635 31.685 119.785 31.835 ;
        RECT 119.635 26.245 119.785 26.395 ;
        RECT 119.635 20.805 119.785 20.955 ;
        RECT 119.635 15.365 119.785 15.515 ;
        RECT 119.635 10.035 119.785 10.185 ;
        RECT 122.395 58.885 122.545 59.035 ;
        RECT 122.395 53.445 122.545 53.595 ;
        RECT 122.395 48.005 122.545 48.155 ;
        RECT 122.395 42.565 122.545 42.715 ;
        RECT 122.395 37.125 122.545 37.275 ;
        RECT 122.395 31.685 122.545 31.835 ;
        RECT 122.395 26.245 122.545 26.395 ;
        RECT 122.395 20.805 122.545 20.955 ;
        RECT 122.395 15.365 122.545 15.515 ;
        RECT 122.395 10.035 122.545 10.185 ;
        RECT 125.155 58.885 125.305 59.035 ;
        RECT 125.155 53.445 125.305 53.595 ;
        RECT 125.155 48.005 125.305 48.155 ;
        RECT 125.155 42.565 125.305 42.715 ;
        RECT 125.155 37.125 125.305 37.275 ;
        RECT 125.155 31.685 125.305 31.835 ;
        RECT 125.155 26.245 125.305 26.395 ;
        RECT 125.155 20.805 125.305 20.955 ;
        RECT 125.155 15.365 125.305 15.515 ;
        RECT 125.155 10.035 125.305 10.185 ;
        RECT 127.915 58.885 128.065 59.035 ;
        RECT 127.915 53.445 128.065 53.595 ;
        RECT 127.915 48.005 128.065 48.155 ;
        RECT 127.915 42.565 128.065 42.715 ;
        RECT 127.915 37.125 128.065 37.275 ;
        RECT 127.915 31.685 128.065 31.835 ;
        RECT 127.915 26.245 128.065 26.395 ;
        RECT 127.915 20.805 128.065 20.955 ;
        RECT 127.915 15.365 128.065 15.515 ;
        RECT 127.915 10.035 128.065 10.185 ;
        RECT 130.675 58.885 130.825 59.035 ;
        RECT 130.675 53.445 130.825 53.595 ;
        RECT 130.675 48.005 130.825 48.155 ;
        RECT 130.675 42.565 130.825 42.715 ;
        RECT 130.675 37.125 130.825 37.275 ;
        RECT 130.675 31.685 130.825 31.835 ;
        RECT 130.675 26.245 130.825 26.395 ;
        RECT 130.675 20.805 130.825 20.955 ;
        RECT 130.675 15.365 130.825 15.515 ;
        RECT 130.675 10.035 130.825 10.185 ;
        RECT 133.435 58.885 133.585 59.035 ;
        RECT 133.435 53.445 133.585 53.595 ;
        RECT 133.435 48.005 133.585 48.155 ;
        RECT 133.435 42.565 133.585 42.715 ;
        RECT 133.435 37.125 133.585 37.275 ;
        RECT 133.435 31.685 133.585 31.835 ;
        RECT 133.435 26.245 133.585 26.395 ;
        RECT 133.435 20.805 133.585 20.955 ;
        RECT 133.435 15.365 133.585 15.515 ;
        RECT 133.435 10.035 133.585 10.185 ;
        RECT 136.195 58.885 136.345 59.035 ;
        RECT 136.195 53.445 136.345 53.595 ;
        RECT 136.195 48.005 136.345 48.155 ;
        RECT 136.195 42.565 136.345 42.715 ;
        RECT 136.195 37.125 136.345 37.275 ;
        RECT 136.195 31.685 136.345 31.835 ;
        RECT 136.195 26.245 136.345 26.395 ;
        RECT 136.195 20.805 136.345 20.955 ;
        RECT 136.195 15.365 136.345 15.515 ;
        RECT 136.195 10.035 136.345 10.185 ;
        RECT 138.955 58.885 139.105 59.035 ;
        RECT 138.955 53.445 139.105 53.595 ;
        RECT 138.955 48.005 139.105 48.155 ;
        RECT 138.955 42.565 139.105 42.715 ;
        RECT 138.955 37.125 139.105 37.275 ;
        RECT 138.955 31.685 139.105 31.835 ;
        RECT 138.955 26.245 139.105 26.395 ;
        RECT 138.955 20.805 139.105 20.955 ;
        RECT 138.955 15.365 139.105 15.515 ;
        RECT 138.955 10.035 139.105 10.185 ;
        RECT 141.715 58.885 141.865 59.035 ;
        RECT 141.715 53.445 141.865 53.595 ;
        RECT 141.715 48.005 141.865 48.155 ;
        RECT 141.715 42.565 141.865 42.715 ;
        RECT 141.715 37.125 141.865 37.275 ;
        RECT 141.715 31.685 141.865 31.835 ;
        RECT 141.715 26.245 141.865 26.395 ;
        RECT 141.715 20.805 141.865 20.955 ;
        RECT 141.715 15.365 141.865 15.515 ;
        RECT 141.715 10.035 141.865 10.185 ;
        RECT 144.475 58.885 144.625 59.035 ;
        RECT 144.475 53.445 144.625 53.595 ;
        RECT 144.475 48.005 144.625 48.155 ;
        RECT 144.475 42.565 144.625 42.715 ;
        RECT 144.475 37.125 144.625 37.275 ;
        RECT 144.475 31.685 144.625 31.835 ;
        RECT 144.475 26.245 144.625 26.395 ;
        RECT 144.475 20.805 144.625 20.955 ;
        RECT 144.475 15.365 144.625 15.515 ;
        RECT 144.475 10.035 144.625 10.185 ;
        RECT 147.235 58.885 147.385 59.035 ;
        RECT 147.235 53.445 147.385 53.595 ;
        RECT 147.235 48.005 147.385 48.155 ;
        RECT 147.235 42.565 147.385 42.715 ;
        RECT 147.235 37.125 147.385 37.275 ;
        RECT 147.235 31.685 147.385 31.835 ;
        RECT 147.235 26.245 147.385 26.395 ;
        RECT 147.235 20.805 147.385 20.955 ;
        RECT 147.235 15.365 147.385 15.515 ;
        RECT 147.235 10.035 147.385 10.185 ;
        RECT 149.995 58.885 150.145 59.035 ;
        RECT 149.995 53.445 150.145 53.595 ;
        RECT 149.995 48.005 150.145 48.155 ;
        RECT 149.995 42.565 150.145 42.715 ;
        RECT 149.995 37.125 150.145 37.275 ;
        RECT 149.995 31.685 150.145 31.835 ;
        RECT 149.995 26.245 150.145 26.395 ;
        RECT 149.995 20.805 150.145 20.955 ;
        RECT 149.995 15.365 150.145 15.515 ;
        RECT 149.995 10.035 150.145 10.185 ;
        RECT 152.755 58.885 152.905 59.035 ;
        RECT 152.755 53.445 152.905 53.595 ;
        RECT 152.755 48.005 152.905 48.155 ;
        RECT 152.755 42.565 152.905 42.715 ;
        RECT 152.755 37.125 152.905 37.275 ;
        RECT 152.755 31.685 152.905 31.835 ;
        RECT 152.755 26.245 152.905 26.395 ;
        RECT 152.755 20.805 152.905 20.955 ;
        RECT 152.755 15.365 152.905 15.515 ;
        RECT 152.755 10.035 152.905 10.185 ;
        RECT 155.515 58.885 155.665 59.035 ;
        RECT 155.515 53.445 155.665 53.595 ;
        RECT 155.515 48.005 155.665 48.155 ;
        RECT 155.515 42.565 155.665 42.715 ;
        RECT 155.515 37.125 155.665 37.275 ;
        RECT 155.515 31.685 155.665 31.835 ;
        RECT 155.515 26.245 155.665 26.395 ;
        RECT 155.515 20.805 155.665 20.955 ;
        RECT 155.515 15.365 155.665 15.515 ;
        RECT 155.515 10.035 155.665 10.185 ;
        RECT 158.275 58.885 158.425 59.035 ;
        RECT 158.275 53.445 158.425 53.595 ;
        RECT 158.275 48.005 158.425 48.155 ;
        RECT 158.275 42.565 158.425 42.715 ;
        RECT 158.275 37.125 158.425 37.275 ;
        RECT 158.275 31.685 158.425 31.835 ;
        RECT 158.275 26.245 158.425 26.395 ;
        RECT 158.275 20.805 158.425 20.955 ;
        RECT 158.275 15.365 158.425 15.515 ;
        RECT 158.275 10.035 158.425 10.185 ;
        RECT 161.035 58.885 161.185 59.035 ;
        RECT 161.035 53.445 161.185 53.595 ;
        RECT 161.035 48.005 161.185 48.155 ;
        RECT 161.035 42.565 161.185 42.715 ;
        RECT 161.035 37.125 161.185 37.275 ;
        RECT 161.035 31.685 161.185 31.835 ;
        RECT 161.035 26.245 161.185 26.395 ;
        RECT 161.035 20.805 161.185 20.955 ;
        RECT 161.035 15.365 161.185 15.515 ;
        RECT 161.035 10.035 161.185 10.185 ;
        RECT 163.795 58.885 163.945 59.035 ;
        RECT 163.795 53.445 163.945 53.595 ;
        RECT 163.795 48.005 163.945 48.155 ;
        RECT 163.795 42.565 163.945 42.715 ;
        RECT 163.795 37.125 163.945 37.275 ;
        RECT 163.795 31.685 163.945 31.835 ;
        RECT 163.795 26.245 163.945 26.395 ;
        RECT 163.795 20.805 163.945 20.955 ;
        RECT 163.795 15.365 163.945 15.515 ;
        RECT 163.795 10.035 163.945 10.185 ;
        RECT 166.555 58.885 166.705 59.035 ;
        RECT 166.555 53.445 166.705 53.595 ;
        RECT 166.555 48.005 166.705 48.155 ;
        RECT 166.555 42.565 166.705 42.715 ;
        RECT 166.555 37.125 166.705 37.275 ;
        RECT 166.555 31.685 166.705 31.835 ;
        RECT 166.555 26.245 166.705 26.395 ;
        RECT 166.555 20.805 166.705 20.955 ;
        RECT 166.555 15.365 166.705 15.515 ;
        RECT 166.555 10.035 166.705 10.185 ;
        RECT 169.315 58.885 169.465 59.035 ;
        RECT 169.315 53.445 169.465 53.595 ;
        RECT 169.315 48.005 169.465 48.155 ;
        RECT 169.315 42.565 169.465 42.715 ;
        RECT 169.315 37.125 169.465 37.275 ;
        RECT 169.315 31.685 169.465 31.835 ;
        RECT 169.315 26.245 169.465 26.395 ;
        RECT 169.315 20.805 169.465 20.955 ;
        RECT 169.315 15.365 169.465 15.515 ;
        RECT 169.315 10.035 169.465 10.185 ;
        RECT 172.075 58.885 172.225 59.035 ;
        RECT 172.075 53.445 172.225 53.595 ;
        RECT 172.075 48.005 172.225 48.155 ;
        RECT 172.075 42.565 172.225 42.715 ;
        RECT 172.075 37.125 172.225 37.275 ;
        RECT 172.075 31.685 172.225 31.835 ;
        RECT 172.075 26.245 172.225 26.395 ;
        RECT 172.075 20.805 172.225 20.955 ;
        RECT 172.075 15.365 172.225 15.515 ;
        RECT 172.075 10.035 172.225 10.185 ;
        RECT 174.835 58.885 174.985 59.035 ;
        RECT 174.835 53.445 174.985 53.595 ;
        RECT 174.835 48.005 174.985 48.155 ;
        RECT 174.835 42.565 174.985 42.715 ;
        RECT 174.835 37.125 174.985 37.275 ;
        RECT 174.835 31.685 174.985 31.835 ;
        RECT 174.835 26.245 174.985 26.395 ;
        RECT 174.835 20.805 174.985 20.955 ;
        RECT 174.835 15.365 174.985 15.515 ;
        RECT 174.835 10.035 174.985 10.185 ;
        RECT 177.595 58.885 177.745 59.035 ;
        RECT 177.595 53.445 177.745 53.595 ;
        RECT 177.595 48.005 177.745 48.155 ;
        RECT 177.595 42.565 177.745 42.715 ;
        RECT 177.595 37.125 177.745 37.275 ;
        RECT 177.595 31.685 177.745 31.835 ;
        RECT 177.595 26.245 177.745 26.395 ;
        RECT 177.595 20.805 177.745 20.955 ;
        RECT 177.595 15.365 177.745 15.515 ;
        RECT 177.595 10.035 177.745 10.185 ;
        RECT 180.355 58.885 180.505 59.035 ;
        RECT 180.355 53.445 180.505 53.595 ;
        RECT 180.355 48.005 180.505 48.155 ;
        RECT 180.355 42.565 180.505 42.715 ;
        RECT 180.355 37.125 180.505 37.275 ;
        RECT 180.355 31.685 180.505 31.835 ;
        RECT 180.355 26.245 180.505 26.395 ;
        RECT 180.355 20.805 180.505 20.955 ;
        RECT 180.355 15.365 180.505 15.515 ;
        RECT 180.355 10.035 180.505 10.185 ;
        RECT 183.115 58.885 183.265 59.035 ;
        RECT 183.115 53.445 183.265 53.595 ;
        RECT 183.115 48.005 183.265 48.155 ;
        RECT 183.115 42.565 183.265 42.715 ;
        RECT 183.115 37.125 183.265 37.275 ;
        RECT 183.115 31.685 183.265 31.835 ;
        RECT 183.115 26.245 183.265 26.395 ;
        RECT 183.115 20.805 183.265 20.955 ;
        RECT 183.115 15.365 183.265 15.515 ;
        RECT 183.115 10.035 183.265 10.185 ;
        RECT 185.875 58.885 186.025 59.035 ;
        RECT 185.875 53.445 186.025 53.595 ;
        RECT 185.875 48.005 186.025 48.155 ;
        RECT 185.875 42.565 186.025 42.715 ;
        RECT 185.875 37.125 186.025 37.275 ;
        RECT 185.875 31.685 186.025 31.835 ;
        RECT 185.875 26.245 186.025 26.395 ;
        RECT 185.875 20.805 186.025 20.955 ;
        RECT 185.875 15.365 186.025 15.515 ;
        RECT 185.875 10.035 186.025 10.185 ;
        RECT 188.635 58.885 188.785 59.035 ;
        RECT 188.635 53.445 188.785 53.595 ;
        RECT 188.635 48.005 188.785 48.155 ;
        RECT 188.635 42.565 188.785 42.715 ;
        RECT 188.635 37.125 188.785 37.275 ;
        RECT 188.635 31.685 188.785 31.835 ;
        RECT 188.635 26.245 188.785 26.395 ;
        RECT 188.635 20.805 188.785 20.955 ;
        RECT 188.635 15.365 188.785 15.515 ;
        RECT 188.635 10.035 188.785 10.185 ;
      LAYER via4 ;
        RECT 13.74 45.3 14.54 46.1 ;
        RECT 13.74 24.9 14.54 25.7 ;
        RECT 19.26 45.3 20.06 46.1 ;
        RECT 19.26 24.9 20.06 25.7 ;
        RECT 24.78 45.3 25.58 46.1 ;
        RECT 24.78 24.9 25.58 25.7 ;
        RECT 30.3 45.3 31.1 46.1 ;
        RECT 30.3 24.9 31.1 25.7 ;
        RECT 35.82 45.3 36.62 46.1 ;
        RECT 35.82 24.9 36.62 25.7 ;
        RECT 41.34 45.3 42.14 46.1 ;
        RECT 41.34 24.9 42.14 25.7 ;
        RECT 46.86 45.3 47.66 46.1 ;
        RECT 46.86 24.9 47.66 25.7 ;
        RECT 52.38 45.3 53.18 46.1 ;
        RECT 52.38 24.9 53.18 25.7 ;
        RECT 57.9 45.3 58.7 46.1 ;
        RECT 57.9 24.9 58.7 25.7 ;
        RECT 63.42 45.3 64.22 46.1 ;
        RECT 63.42 24.9 64.22 25.7 ;
        RECT 68.94 45.3 69.74 46.1 ;
        RECT 68.94 24.9 69.74 25.7 ;
        RECT 74.46 45.3 75.26 46.1 ;
        RECT 74.46 24.9 75.26 25.7 ;
        RECT 79.98 45.3 80.78 46.1 ;
        RECT 79.98 24.9 80.78 25.7 ;
        RECT 85.5 45.3 86.3 46.1 ;
        RECT 85.5 24.9 86.3 25.7 ;
        RECT 91.02 45.3 91.82 46.1 ;
        RECT 91.02 24.9 91.82 25.7 ;
        RECT 96.54 45.3 97.34 46.1 ;
        RECT 96.54 24.9 97.34 25.7 ;
        RECT 102.06 45.3 102.86 46.1 ;
        RECT 102.06 24.9 102.86 25.7 ;
        RECT 107.58 45.3 108.38 46.1 ;
        RECT 107.58 24.9 108.38 25.7 ;
        RECT 113.1 45.3 113.9 46.1 ;
        RECT 113.1 24.9 113.9 25.7 ;
        RECT 118.62 45.3 119.42 46.1 ;
        RECT 118.62 24.9 119.42 25.7 ;
        RECT 124.14 45.3 124.94 46.1 ;
        RECT 124.14 24.9 124.94 25.7 ;
        RECT 129.66 45.3 130.46 46.1 ;
        RECT 129.66 24.9 130.46 25.7 ;
        RECT 135.18 45.3 135.98 46.1 ;
        RECT 135.18 24.9 135.98 25.7 ;
        RECT 140.7 45.3 141.5 46.1 ;
        RECT 140.7 24.9 141.5 25.7 ;
        RECT 146.22 45.3 147.02 46.1 ;
        RECT 146.22 24.9 147.02 25.7 ;
        RECT 151.74 45.3 152.54 46.1 ;
        RECT 151.74 24.9 152.54 25.7 ;
        RECT 157.26 45.3 158.06 46.1 ;
        RECT 157.26 24.9 158.06 25.7 ;
        RECT 162.78 45.3 163.58 46.1 ;
        RECT 162.78 24.9 163.58 25.7 ;
        RECT 168.3 45.3 169.1 46.1 ;
        RECT 168.3 24.9 169.1 25.7 ;
        RECT 173.82 45.3 174.62 46.1 ;
        RECT 173.82 24.9 174.62 25.7 ;
        RECT 179.34 45.3 180.14 46.1 ;
        RECT 179.34 24.9 180.14 25.7 ;
        RECT 184.86 45.3 185.66 46.1 ;
        RECT 184.86 24.9 185.66 25.7 ;
      LAYER mcon ;
        RECT 148.145 58.875 148.315 59.045 ;
        RECT 148.145 53.435 148.315 53.605 ;
        RECT 148.145 47.995 148.315 48.165 ;
        RECT 148.145 42.555 148.315 42.725 ;
        RECT 148.145 37.115 148.315 37.285 ;
        RECT 148.145 31.675 148.315 31.845 ;
        RECT 148.145 26.235 148.315 26.405 ;
        RECT 148.145 20.795 148.315 20.965 ;
        RECT 148.145 15.355 148.315 15.525 ;
        RECT 148.145 9.915 148.315 10.085 ;
        RECT 148.605 58.875 148.775 59.045 ;
        RECT 148.605 53.435 148.775 53.605 ;
        RECT 148.605 47.995 148.775 48.165 ;
        RECT 148.605 42.555 148.775 42.725 ;
        RECT 148.605 37.115 148.775 37.285 ;
        RECT 148.605 31.675 148.775 31.845 ;
        RECT 148.605 26.235 148.775 26.405 ;
        RECT 148.605 20.795 148.775 20.965 ;
        RECT 148.605 15.355 148.775 15.525 ;
        RECT 148.605 9.915 148.775 10.085 ;
        RECT 149.065 58.875 149.235 59.045 ;
        RECT 149.065 53.435 149.235 53.605 ;
        RECT 149.065 47.995 149.235 48.165 ;
        RECT 149.065 42.555 149.235 42.725 ;
        RECT 149.065 37.115 149.235 37.285 ;
        RECT 149.065 31.675 149.235 31.845 ;
        RECT 149.065 26.235 149.235 26.405 ;
        RECT 149.065 20.795 149.235 20.965 ;
        RECT 149.065 15.355 149.235 15.525 ;
        RECT 149.065 9.915 149.235 10.085 ;
        RECT 149.525 58.875 149.695 59.045 ;
        RECT 149.525 53.435 149.695 53.605 ;
        RECT 149.525 47.995 149.695 48.165 ;
        RECT 149.525 42.555 149.695 42.725 ;
        RECT 149.525 37.115 149.695 37.285 ;
        RECT 149.525 31.675 149.695 31.845 ;
        RECT 149.525 26.235 149.695 26.405 ;
        RECT 149.525 20.795 149.695 20.965 ;
        RECT 149.525 15.355 149.695 15.525 ;
        RECT 149.525 9.915 149.695 10.085 ;
        RECT 149.985 58.875 150.155 59.045 ;
        RECT 149.985 53.435 150.155 53.605 ;
        RECT 149.985 47.995 150.155 48.165 ;
        RECT 149.985 42.555 150.155 42.725 ;
        RECT 149.985 37.115 150.155 37.285 ;
        RECT 149.985 31.675 150.155 31.845 ;
        RECT 149.985 26.235 150.155 26.405 ;
        RECT 149.985 20.795 150.155 20.965 ;
        RECT 149.985 15.355 150.155 15.525 ;
        RECT 149.985 9.915 150.155 10.085 ;
        RECT 150.445 58.875 150.615 59.045 ;
        RECT 150.445 53.435 150.615 53.605 ;
        RECT 150.445 47.995 150.615 48.165 ;
        RECT 150.445 42.555 150.615 42.725 ;
        RECT 150.445 37.115 150.615 37.285 ;
        RECT 150.445 31.675 150.615 31.845 ;
        RECT 150.445 26.235 150.615 26.405 ;
        RECT 150.445 20.795 150.615 20.965 ;
        RECT 150.445 15.355 150.615 15.525 ;
        RECT 150.445 9.915 150.615 10.085 ;
        RECT 150.905 58.875 151.075 59.045 ;
        RECT 150.905 53.435 151.075 53.605 ;
        RECT 150.905 47.995 151.075 48.165 ;
        RECT 150.905 42.555 151.075 42.725 ;
        RECT 150.905 37.115 151.075 37.285 ;
        RECT 150.905 31.675 151.075 31.845 ;
        RECT 150.905 26.235 151.075 26.405 ;
        RECT 150.905 20.795 151.075 20.965 ;
        RECT 150.905 15.355 151.075 15.525 ;
        RECT 150.905 9.915 151.075 10.085 ;
        RECT 151.365 58.875 151.535 59.045 ;
        RECT 151.365 53.435 151.535 53.605 ;
        RECT 151.365 47.995 151.535 48.165 ;
        RECT 151.365 42.555 151.535 42.725 ;
        RECT 151.365 37.115 151.535 37.285 ;
        RECT 151.365 31.675 151.535 31.845 ;
        RECT 151.365 26.235 151.535 26.405 ;
        RECT 151.365 20.795 151.535 20.965 ;
        RECT 151.365 15.355 151.535 15.525 ;
        RECT 151.365 9.915 151.535 10.085 ;
        RECT 151.825 58.875 151.995 59.045 ;
        RECT 151.825 53.435 151.995 53.605 ;
        RECT 151.825 47.995 151.995 48.165 ;
        RECT 151.825 42.555 151.995 42.725 ;
        RECT 151.825 37.115 151.995 37.285 ;
        RECT 151.825 31.675 151.995 31.845 ;
        RECT 151.825 26.235 151.995 26.405 ;
        RECT 151.825 20.795 151.995 20.965 ;
        RECT 151.825 15.355 151.995 15.525 ;
        RECT 151.825 9.915 151.995 10.085 ;
        RECT 152.285 58.875 152.455 59.045 ;
        RECT 152.285 53.435 152.455 53.605 ;
        RECT 152.285 47.995 152.455 48.165 ;
        RECT 152.285 42.555 152.455 42.725 ;
        RECT 152.285 37.115 152.455 37.285 ;
        RECT 152.285 31.675 152.455 31.845 ;
        RECT 152.285 26.235 152.455 26.405 ;
        RECT 152.285 20.795 152.455 20.965 ;
        RECT 152.285 15.355 152.455 15.525 ;
        RECT 152.285 9.915 152.455 10.085 ;
        RECT 152.745 58.875 152.915 59.045 ;
        RECT 152.745 53.435 152.915 53.605 ;
        RECT 152.745 47.995 152.915 48.165 ;
        RECT 152.745 42.555 152.915 42.725 ;
        RECT 152.745 37.115 152.915 37.285 ;
        RECT 152.745 31.675 152.915 31.845 ;
        RECT 152.745 26.235 152.915 26.405 ;
        RECT 152.745 20.795 152.915 20.965 ;
        RECT 152.745 15.355 152.915 15.525 ;
        RECT 152.745 9.915 152.915 10.085 ;
        RECT 153.205 58.875 153.375 59.045 ;
        RECT 153.205 53.435 153.375 53.605 ;
        RECT 153.205 47.995 153.375 48.165 ;
        RECT 153.205 42.555 153.375 42.725 ;
        RECT 153.205 37.115 153.375 37.285 ;
        RECT 153.205 31.675 153.375 31.845 ;
        RECT 153.205 26.235 153.375 26.405 ;
        RECT 153.205 20.795 153.375 20.965 ;
        RECT 153.205 15.355 153.375 15.525 ;
        RECT 153.205 9.915 153.375 10.085 ;
        RECT 153.665 58.875 153.835 59.045 ;
        RECT 153.665 53.435 153.835 53.605 ;
        RECT 153.665 47.995 153.835 48.165 ;
        RECT 153.665 42.555 153.835 42.725 ;
        RECT 153.665 37.115 153.835 37.285 ;
        RECT 153.665 31.675 153.835 31.845 ;
        RECT 153.665 26.235 153.835 26.405 ;
        RECT 153.665 20.795 153.835 20.965 ;
        RECT 153.665 15.355 153.835 15.525 ;
        RECT 153.665 9.915 153.835 10.085 ;
        RECT 154.125 58.875 154.295 59.045 ;
        RECT 154.125 53.435 154.295 53.605 ;
        RECT 154.125 47.995 154.295 48.165 ;
        RECT 154.125 42.555 154.295 42.725 ;
        RECT 154.125 37.115 154.295 37.285 ;
        RECT 154.125 31.675 154.295 31.845 ;
        RECT 154.125 26.235 154.295 26.405 ;
        RECT 154.125 20.795 154.295 20.965 ;
        RECT 154.125 15.355 154.295 15.525 ;
        RECT 154.125 9.915 154.295 10.085 ;
        RECT 154.585 58.875 154.755 59.045 ;
        RECT 154.585 53.435 154.755 53.605 ;
        RECT 154.585 47.995 154.755 48.165 ;
        RECT 154.585 42.555 154.755 42.725 ;
        RECT 154.585 37.115 154.755 37.285 ;
        RECT 154.585 31.675 154.755 31.845 ;
        RECT 154.585 26.235 154.755 26.405 ;
        RECT 154.585 20.795 154.755 20.965 ;
        RECT 154.585 15.355 154.755 15.525 ;
        RECT 154.585 9.915 154.755 10.085 ;
        RECT 155.045 58.875 155.215 59.045 ;
        RECT 155.045 53.435 155.215 53.605 ;
        RECT 155.045 47.995 155.215 48.165 ;
        RECT 155.045 42.555 155.215 42.725 ;
        RECT 155.045 37.115 155.215 37.285 ;
        RECT 155.045 31.675 155.215 31.845 ;
        RECT 155.045 26.235 155.215 26.405 ;
        RECT 155.045 20.795 155.215 20.965 ;
        RECT 155.045 15.355 155.215 15.525 ;
        RECT 155.045 9.915 155.215 10.085 ;
        RECT 155.505 58.875 155.675 59.045 ;
        RECT 155.505 53.435 155.675 53.605 ;
        RECT 155.505 47.995 155.675 48.165 ;
        RECT 155.505 42.555 155.675 42.725 ;
        RECT 155.505 37.115 155.675 37.285 ;
        RECT 155.505 31.675 155.675 31.845 ;
        RECT 155.505 26.235 155.675 26.405 ;
        RECT 155.505 20.795 155.675 20.965 ;
        RECT 155.505 15.355 155.675 15.525 ;
        RECT 155.505 9.915 155.675 10.085 ;
        RECT 155.965 58.875 156.135 59.045 ;
        RECT 155.965 53.435 156.135 53.605 ;
        RECT 155.965 47.995 156.135 48.165 ;
        RECT 155.965 42.555 156.135 42.725 ;
        RECT 155.965 37.115 156.135 37.285 ;
        RECT 155.965 31.675 156.135 31.845 ;
        RECT 155.965 26.235 156.135 26.405 ;
        RECT 155.965 20.795 156.135 20.965 ;
        RECT 155.965 15.355 156.135 15.525 ;
        RECT 155.965 9.915 156.135 10.085 ;
        RECT 156.425 58.875 156.595 59.045 ;
        RECT 156.425 53.435 156.595 53.605 ;
        RECT 156.425 47.995 156.595 48.165 ;
        RECT 156.425 42.555 156.595 42.725 ;
        RECT 156.425 37.115 156.595 37.285 ;
        RECT 156.425 31.675 156.595 31.845 ;
        RECT 156.425 26.235 156.595 26.405 ;
        RECT 156.425 20.795 156.595 20.965 ;
        RECT 156.425 15.355 156.595 15.525 ;
        RECT 156.425 9.915 156.595 10.085 ;
        RECT 156.885 58.875 157.055 59.045 ;
        RECT 156.885 53.435 157.055 53.605 ;
        RECT 156.885 47.995 157.055 48.165 ;
        RECT 156.885 42.555 157.055 42.725 ;
        RECT 156.885 37.115 157.055 37.285 ;
        RECT 156.885 31.675 157.055 31.845 ;
        RECT 156.885 26.235 157.055 26.405 ;
        RECT 156.885 20.795 157.055 20.965 ;
        RECT 156.885 15.355 157.055 15.525 ;
        RECT 156.885 9.915 157.055 10.085 ;
        RECT 157.345 58.875 157.515 59.045 ;
        RECT 157.345 53.435 157.515 53.605 ;
        RECT 157.345 47.995 157.515 48.165 ;
        RECT 157.345 42.555 157.515 42.725 ;
        RECT 157.345 37.115 157.515 37.285 ;
        RECT 157.345 31.675 157.515 31.845 ;
        RECT 157.345 26.235 157.515 26.405 ;
        RECT 157.345 20.795 157.515 20.965 ;
        RECT 157.345 15.355 157.515 15.525 ;
        RECT 157.345 9.915 157.515 10.085 ;
        RECT 157.805 58.875 157.975 59.045 ;
        RECT 157.805 53.435 157.975 53.605 ;
        RECT 157.805 47.995 157.975 48.165 ;
        RECT 157.805 42.555 157.975 42.725 ;
        RECT 157.805 37.115 157.975 37.285 ;
        RECT 157.805 31.675 157.975 31.845 ;
        RECT 157.805 26.235 157.975 26.405 ;
        RECT 157.805 20.795 157.975 20.965 ;
        RECT 157.805 15.355 157.975 15.525 ;
        RECT 157.805 9.915 157.975 10.085 ;
        RECT 158.265 58.875 158.435 59.045 ;
        RECT 158.265 53.435 158.435 53.605 ;
        RECT 158.265 47.995 158.435 48.165 ;
        RECT 158.265 42.555 158.435 42.725 ;
        RECT 158.265 37.115 158.435 37.285 ;
        RECT 158.265 31.675 158.435 31.845 ;
        RECT 158.265 26.235 158.435 26.405 ;
        RECT 158.265 20.795 158.435 20.965 ;
        RECT 158.265 15.355 158.435 15.525 ;
        RECT 158.265 9.915 158.435 10.085 ;
        RECT 158.725 58.875 158.895 59.045 ;
        RECT 158.725 53.435 158.895 53.605 ;
        RECT 158.725 47.995 158.895 48.165 ;
        RECT 158.725 42.555 158.895 42.725 ;
        RECT 158.725 37.115 158.895 37.285 ;
        RECT 158.725 31.675 158.895 31.845 ;
        RECT 158.725 26.235 158.895 26.405 ;
        RECT 158.725 20.795 158.895 20.965 ;
        RECT 158.725 15.355 158.895 15.525 ;
        RECT 158.725 9.915 158.895 10.085 ;
        RECT 159.185 58.875 159.355 59.045 ;
        RECT 159.185 53.435 159.355 53.605 ;
        RECT 159.185 47.995 159.355 48.165 ;
        RECT 159.185 42.555 159.355 42.725 ;
        RECT 159.185 37.115 159.355 37.285 ;
        RECT 159.185 31.675 159.355 31.845 ;
        RECT 159.185 26.235 159.355 26.405 ;
        RECT 159.185 20.795 159.355 20.965 ;
        RECT 159.185 15.355 159.355 15.525 ;
        RECT 159.185 9.915 159.355 10.085 ;
        RECT 159.645 58.875 159.815 59.045 ;
        RECT 159.645 53.435 159.815 53.605 ;
        RECT 159.645 47.995 159.815 48.165 ;
        RECT 159.645 42.555 159.815 42.725 ;
        RECT 159.645 37.115 159.815 37.285 ;
        RECT 159.645 31.675 159.815 31.845 ;
        RECT 159.645 26.235 159.815 26.405 ;
        RECT 159.645 20.795 159.815 20.965 ;
        RECT 159.645 15.355 159.815 15.525 ;
        RECT 159.645 9.915 159.815 10.085 ;
        RECT 160.105 58.875 160.275 59.045 ;
        RECT 160.105 53.435 160.275 53.605 ;
        RECT 160.105 47.995 160.275 48.165 ;
        RECT 160.105 42.555 160.275 42.725 ;
        RECT 160.105 37.115 160.275 37.285 ;
        RECT 160.105 31.675 160.275 31.845 ;
        RECT 160.105 26.235 160.275 26.405 ;
        RECT 160.105 20.795 160.275 20.965 ;
        RECT 160.105 15.355 160.275 15.525 ;
        RECT 160.105 9.915 160.275 10.085 ;
        RECT 160.565 58.875 160.735 59.045 ;
        RECT 160.565 53.435 160.735 53.605 ;
        RECT 160.565 47.995 160.735 48.165 ;
        RECT 160.565 42.555 160.735 42.725 ;
        RECT 160.565 37.115 160.735 37.285 ;
        RECT 160.565 31.675 160.735 31.845 ;
        RECT 160.565 26.235 160.735 26.405 ;
        RECT 160.565 20.795 160.735 20.965 ;
        RECT 160.565 15.355 160.735 15.525 ;
        RECT 160.565 9.915 160.735 10.085 ;
        RECT 161.025 58.875 161.195 59.045 ;
        RECT 161.025 53.435 161.195 53.605 ;
        RECT 161.025 47.995 161.195 48.165 ;
        RECT 161.025 42.555 161.195 42.725 ;
        RECT 161.025 37.115 161.195 37.285 ;
        RECT 161.025 31.675 161.195 31.845 ;
        RECT 161.025 26.235 161.195 26.405 ;
        RECT 161.025 20.795 161.195 20.965 ;
        RECT 161.025 15.355 161.195 15.525 ;
        RECT 161.025 9.915 161.195 10.085 ;
        RECT 161.485 58.875 161.655 59.045 ;
        RECT 161.485 53.435 161.655 53.605 ;
        RECT 161.485 47.995 161.655 48.165 ;
        RECT 161.485 42.555 161.655 42.725 ;
        RECT 161.485 37.115 161.655 37.285 ;
        RECT 161.485 31.675 161.655 31.845 ;
        RECT 161.485 26.235 161.655 26.405 ;
        RECT 161.485 20.795 161.655 20.965 ;
        RECT 161.485 15.355 161.655 15.525 ;
        RECT 161.485 9.915 161.655 10.085 ;
        RECT 161.945 58.875 162.115 59.045 ;
        RECT 161.945 53.435 162.115 53.605 ;
        RECT 161.945 47.995 162.115 48.165 ;
        RECT 161.945 42.555 162.115 42.725 ;
        RECT 161.945 37.115 162.115 37.285 ;
        RECT 161.945 31.675 162.115 31.845 ;
        RECT 161.945 26.235 162.115 26.405 ;
        RECT 161.945 20.795 162.115 20.965 ;
        RECT 161.945 15.355 162.115 15.525 ;
        RECT 161.945 9.915 162.115 10.085 ;
        RECT 162.405 58.875 162.575 59.045 ;
        RECT 162.405 53.435 162.575 53.605 ;
        RECT 162.405 47.995 162.575 48.165 ;
        RECT 162.405 42.555 162.575 42.725 ;
        RECT 162.405 37.115 162.575 37.285 ;
        RECT 162.405 31.675 162.575 31.845 ;
        RECT 162.405 26.235 162.575 26.405 ;
        RECT 162.405 20.795 162.575 20.965 ;
        RECT 162.405 15.355 162.575 15.525 ;
        RECT 162.405 9.915 162.575 10.085 ;
        RECT 162.865 58.875 163.035 59.045 ;
        RECT 162.865 53.435 163.035 53.605 ;
        RECT 162.865 47.995 163.035 48.165 ;
        RECT 162.865 42.555 163.035 42.725 ;
        RECT 162.865 37.115 163.035 37.285 ;
        RECT 162.865 31.675 163.035 31.845 ;
        RECT 162.865 26.235 163.035 26.405 ;
        RECT 162.865 20.795 163.035 20.965 ;
        RECT 162.865 15.355 163.035 15.525 ;
        RECT 162.865 9.915 163.035 10.085 ;
        RECT 163.325 58.875 163.495 59.045 ;
        RECT 163.325 53.435 163.495 53.605 ;
        RECT 163.325 47.995 163.495 48.165 ;
        RECT 163.325 42.555 163.495 42.725 ;
        RECT 163.325 37.115 163.495 37.285 ;
        RECT 163.325 31.675 163.495 31.845 ;
        RECT 163.325 26.235 163.495 26.405 ;
        RECT 163.325 20.795 163.495 20.965 ;
        RECT 163.325 15.355 163.495 15.525 ;
        RECT 163.325 9.915 163.495 10.085 ;
        RECT 163.785 58.875 163.955 59.045 ;
        RECT 163.785 53.435 163.955 53.605 ;
        RECT 163.785 47.995 163.955 48.165 ;
        RECT 163.785 42.555 163.955 42.725 ;
        RECT 163.785 37.115 163.955 37.285 ;
        RECT 163.785 31.675 163.955 31.845 ;
        RECT 163.785 26.235 163.955 26.405 ;
        RECT 163.785 20.795 163.955 20.965 ;
        RECT 163.785 15.355 163.955 15.525 ;
        RECT 163.785 9.915 163.955 10.085 ;
        RECT 164.245 58.875 164.415 59.045 ;
        RECT 164.245 53.435 164.415 53.605 ;
        RECT 164.245 47.995 164.415 48.165 ;
        RECT 164.245 42.555 164.415 42.725 ;
        RECT 164.245 37.115 164.415 37.285 ;
        RECT 164.245 31.675 164.415 31.845 ;
        RECT 164.245 26.235 164.415 26.405 ;
        RECT 164.245 20.795 164.415 20.965 ;
        RECT 164.245 15.355 164.415 15.525 ;
        RECT 164.245 9.915 164.415 10.085 ;
        RECT 164.705 58.875 164.875 59.045 ;
        RECT 164.705 53.435 164.875 53.605 ;
        RECT 164.705 47.995 164.875 48.165 ;
        RECT 164.705 42.555 164.875 42.725 ;
        RECT 164.705 37.115 164.875 37.285 ;
        RECT 164.705 31.675 164.875 31.845 ;
        RECT 164.705 26.235 164.875 26.405 ;
        RECT 164.705 20.795 164.875 20.965 ;
        RECT 164.705 15.355 164.875 15.525 ;
        RECT 164.705 9.915 164.875 10.085 ;
        RECT 165.165 58.875 165.335 59.045 ;
        RECT 165.165 53.435 165.335 53.605 ;
        RECT 165.165 47.995 165.335 48.165 ;
        RECT 165.165 42.555 165.335 42.725 ;
        RECT 165.165 37.115 165.335 37.285 ;
        RECT 165.165 31.675 165.335 31.845 ;
        RECT 165.165 26.235 165.335 26.405 ;
        RECT 165.165 20.795 165.335 20.965 ;
        RECT 165.165 15.355 165.335 15.525 ;
        RECT 165.165 9.915 165.335 10.085 ;
        RECT 165.625 58.875 165.795 59.045 ;
        RECT 165.625 53.435 165.795 53.605 ;
        RECT 165.625 47.995 165.795 48.165 ;
        RECT 165.625 42.555 165.795 42.725 ;
        RECT 165.625 37.115 165.795 37.285 ;
        RECT 165.625 31.675 165.795 31.845 ;
        RECT 165.625 26.235 165.795 26.405 ;
        RECT 165.625 20.795 165.795 20.965 ;
        RECT 165.625 15.355 165.795 15.525 ;
        RECT 165.625 9.915 165.795 10.085 ;
        RECT 166.085 58.875 166.255 59.045 ;
        RECT 166.085 53.435 166.255 53.605 ;
        RECT 166.085 47.995 166.255 48.165 ;
        RECT 166.085 42.555 166.255 42.725 ;
        RECT 166.085 37.115 166.255 37.285 ;
        RECT 166.085 31.675 166.255 31.845 ;
        RECT 166.085 26.235 166.255 26.405 ;
        RECT 166.085 20.795 166.255 20.965 ;
        RECT 166.085 15.355 166.255 15.525 ;
        RECT 166.085 9.915 166.255 10.085 ;
        RECT 166.545 58.875 166.715 59.045 ;
        RECT 166.545 53.435 166.715 53.605 ;
        RECT 166.545 47.995 166.715 48.165 ;
        RECT 166.545 42.555 166.715 42.725 ;
        RECT 166.545 37.115 166.715 37.285 ;
        RECT 166.545 31.675 166.715 31.845 ;
        RECT 166.545 26.235 166.715 26.405 ;
        RECT 166.545 20.795 166.715 20.965 ;
        RECT 166.545 15.355 166.715 15.525 ;
        RECT 166.545 9.915 166.715 10.085 ;
        RECT 167.005 58.875 167.175 59.045 ;
        RECT 167.005 53.435 167.175 53.605 ;
        RECT 167.005 47.995 167.175 48.165 ;
        RECT 167.005 42.555 167.175 42.725 ;
        RECT 167.005 37.115 167.175 37.285 ;
        RECT 167.005 31.675 167.175 31.845 ;
        RECT 167.005 26.235 167.175 26.405 ;
        RECT 167.005 20.795 167.175 20.965 ;
        RECT 167.005 15.355 167.175 15.525 ;
        RECT 167.005 9.915 167.175 10.085 ;
        RECT 167.465 58.875 167.635 59.045 ;
        RECT 167.465 53.435 167.635 53.605 ;
        RECT 167.465 47.995 167.635 48.165 ;
        RECT 167.465 42.555 167.635 42.725 ;
        RECT 167.465 37.115 167.635 37.285 ;
        RECT 167.465 31.675 167.635 31.845 ;
        RECT 167.465 26.235 167.635 26.405 ;
        RECT 167.465 20.795 167.635 20.965 ;
        RECT 167.465 15.355 167.635 15.525 ;
        RECT 167.465 9.915 167.635 10.085 ;
        RECT 167.925 58.875 168.095 59.045 ;
        RECT 167.925 53.435 168.095 53.605 ;
        RECT 167.925 47.995 168.095 48.165 ;
        RECT 167.925 42.555 168.095 42.725 ;
        RECT 167.925 37.115 168.095 37.285 ;
        RECT 167.925 31.675 168.095 31.845 ;
        RECT 167.925 26.235 168.095 26.405 ;
        RECT 167.925 20.795 168.095 20.965 ;
        RECT 167.925 15.355 168.095 15.525 ;
        RECT 167.925 9.915 168.095 10.085 ;
        RECT 168.385 58.875 168.555 59.045 ;
        RECT 168.385 53.435 168.555 53.605 ;
        RECT 168.385 47.995 168.555 48.165 ;
        RECT 168.385 42.555 168.555 42.725 ;
        RECT 168.385 37.115 168.555 37.285 ;
        RECT 168.385 31.675 168.555 31.845 ;
        RECT 168.385 26.235 168.555 26.405 ;
        RECT 168.385 20.795 168.555 20.965 ;
        RECT 168.385 15.355 168.555 15.525 ;
        RECT 168.385 9.915 168.555 10.085 ;
        RECT 168.845 58.875 169.015 59.045 ;
        RECT 168.845 53.435 169.015 53.605 ;
        RECT 168.845 47.995 169.015 48.165 ;
        RECT 168.845 42.555 169.015 42.725 ;
        RECT 168.845 37.115 169.015 37.285 ;
        RECT 168.845 31.675 169.015 31.845 ;
        RECT 168.845 26.235 169.015 26.405 ;
        RECT 168.845 20.795 169.015 20.965 ;
        RECT 168.845 15.355 169.015 15.525 ;
        RECT 168.845 9.915 169.015 10.085 ;
        RECT 169.305 58.875 169.475 59.045 ;
        RECT 169.305 53.435 169.475 53.605 ;
        RECT 169.305 47.995 169.475 48.165 ;
        RECT 169.305 42.555 169.475 42.725 ;
        RECT 169.305 37.115 169.475 37.285 ;
        RECT 169.305 31.675 169.475 31.845 ;
        RECT 169.305 26.235 169.475 26.405 ;
        RECT 169.305 20.795 169.475 20.965 ;
        RECT 169.305 15.355 169.475 15.525 ;
        RECT 169.305 9.915 169.475 10.085 ;
        RECT 169.765 58.875 169.935 59.045 ;
        RECT 169.765 53.435 169.935 53.605 ;
        RECT 169.765 47.995 169.935 48.165 ;
        RECT 169.765 42.555 169.935 42.725 ;
        RECT 169.765 37.115 169.935 37.285 ;
        RECT 169.765 31.675 169.935 31.845 ;
        RECT 169.765 26.235 169.935 26.405 ;
        RECT 169.765 20.795 169.935 20.965 ;
        RECT 169.765 15.355 169.935 15.525 ;
        RECT 169.765 9.915 169.935 10.085 ;
        RECT 170.225 58.875 170.395 59.045 ;
        RECT 170.225 53.435 170.395 53.605 ;
        RECT 170.225 47.995 170.395 48.165 ;
        RECT 170.225 42.555 170.395 42.725 ;
        RECT 170.225 37.115 170.395 37.285 ;
        RECT 170.225 31.675 170.395 31.845 ;
        RECT 170.225 26.235 170.395 26.405 ;
        RECT 170.225 20.795 170.395 20.965 ;
        RECT 170.225 15.355 170.395 15.525 ;
        RECT 170.225 9.915 170.395 10.085 ;
        RECT 170.685 58.875 170.855 59.045 ;
        RECT 170.685 53.435 170.855 53.605 ;
        RECT 170.685 47.995 170.855 48.165 ;
        RECT 170.685 42.555 170.855 42.725 ;
        RECT 170.685 37.115 170.855 37.285 ;
        RECT 170.685 31.675 170.855 31.845 ;
        RECT 170.685 26.235 170.855 26.405 ;
        RECT 170.685 20.795 170.855 20.965 ;
        RECT 170.685 15.355 170.855 15.525 ;
        RECT 170.685 9.915 170.855 10.085 ;
        RECT 171.145 58.875 171.315 59.045 ;
        RECT 171.145 53.435 171.315 53.605 ;
        RECT 171.145 47.995 171.315 48.165 ;
        RECT 171.145 42.555 171.315 42.725 ;
        RECT 171.145 37.115 171.315 37.285 ;
        RECT 171.145 31.675 171.315 31.845 ;
        RECT 171.145 26.235 171.315 26.405 ;
        RECT 171.145 20.795 171.315 20.965 ;
        RECT 171.145 15.355 171.315 15.525 ;
        RECT 171.145 9.915 171.315 10.085 ;
        RECT 171.605 58.875 171.775 59.045 ;
        RECT 171.605 53.435 171.775 53.605 ;
        RECT 171.605 47.995 171.775 48.165 ;
        RECT 171.605 42.555 171.775 42.725 ;
        RECT 171.605 37.115 171.775 37.285 ;
        RECT 171.605 31.675 171.775 31.845 ;
        RECT 171.605 26.235 171.775 26.405 ;
        RECT 171.605 20.795 171.775 20.965 ;
        RECT 171.605 15.355 171.775 15.525 ;
        RECT 171.605 9.915 171.775 10.085 ;
        RECT 172.065 58.875 172.235 59.045 ;
        RECT 172.065 53.435 172.235 53.605 ;
        RECT 172.065 47.995 172.235 48.165 ;
        RECT 172.065 42.555 172.235 42.725 ;
        RECT 172.065 37.115 172.235 37.285 ;
        RECT 172.065 31.675 172.235 31.845 ;
        RECT 172.065 26.235 172.235 26.405 ;
        RECT 172.065 20.795 172.235 20.965 ;
        RECT 172.065 15.355 172.235 15.525 ;
        RECT 172.065 9.915 172.235 10.085 ;
        RECT 172.525 58.875 172.695 59.045 ;
        RECT 172.525 53.435 172.695 53.605 ;
        RECT 172.525 47.995 172.695 48.165 ;
        RECT 172.525 42.555 172.695 42.725 ;
        RECT 172.525 37.115 172.695 37.285 ;
        RECT 172.525 31.675 172.695 31.845 ;
        RECT 172.525 26.235 172.695 26.405 ;
        RECT 172.525 20.795 172.695 20.965 ;
        RECT 172.525 15.355 172.695 15.525 ;
        RECT 172.525 9.915 172.695 10.085 ;
        RECT 172.985 58.875 173.155 59.045 ;
        RECT 172.985 53.435 173.155 53.605 ;
        RECT 172.985 47.995 173.155 48.165 ;
        RECT 172.985 42.555 173.155 42.725 ;
        RECT 172.985 37.115 173.155 37.285 ;
        RECT 172.985 31.675 173.155 31.845 ;
        RECT 172.985 26.235 173.155 26.405 ;
        RECT 172.985 20.795 173.155 20.965 ;
        RECT 172.985 15.355 173.155 15.525 ;
        RECT 172.985 9.915 173.155 10.085 ;
        RECT 173.445 58.875 173.615 59.045 ;
        RECT 173.445 53.435 173.615 53.605 ;
        RECT 173.445 47.995 173.615 48.165 ;
        RECT 173.445 42.555 173.615 42.725 ;
        RECT 173.445 37.115 173.615 37.285 ;
        RECT 173.445 31.675 173.615 31.845 ;
        RECT 173.445 26.235 173.615 26.405 ;
        RECT 173.445 20.795 173.615 20.965 ;
        RECT 173.445 15.355 173.615 15.525 ;
        RECT 173.445 9.915 173.615 10.085 ;
        RECT 173.905 58.875 174.075 59.045 ;
        RECT 173.905 53.435 174.075 53.605 ;
        RECT 173.905 47.995 174.075 48.165 ;
        RECT 173.905 42.555 174.075 42.725 ;
        RECT 173.905 37.115 174.075 37.285 ;
        RECT 173.905 31.675 174.075 31.845 ;
        RECT 173.905 26.235 174.075 26.405 ;
        RECT 173.905 20.795 174.075 20.965 ;
        RECT 173.905 15.355 174.075 15.525 ;
        RECT 173.905 9.915 174.075 10.085 ;
        RECT 174.365 58.875 174.535 59.045 ;
        RECT 174.365 53.435 174.535 53.605 ;
        RECT 174.365 47.995 174.535 48.165 ;
        RECT 174.365 42.555 174.535 42.725 ;
        RECT 174.365 37.115 174.535 37.285 ;
        RECT 174.365 31.675 174.535 31.845 ;
        RECT 174.365 26.235 174.535 26.405 ;
        RECT 174.365 20.795 174.535 20.965 ;
        RECT 174.365 15.355 174.535 15.525 ;
        RECT 174.365 9.915 174.535 10.085 ;
        RECT 174.825 58.875 174.995 59.045 ;
        RECT 174.825 53.435 174.995 53.605 ;
        RECT 174.825 47.995 174.995 48.165 ;
        RECT 174.825 42.555 174.995 42.725 ;
        RECT 174.825 37.115 174.995 37.285 ;
        RECT 174.825 31.675 174.995 31.845 ;
        RECT 174.825 26.235 174.995 26.405 ;
        RECT 174.825 20.795 174.995 20.965 ;
        RECT 174.825 15.355 174.995 15.525 ;
        RECT 174.825 9.915 174.995 10.085 ;
        RECT 175.285 58.875 175.455 59.045 ;
        RECT 175.285 53.435 175.455 53.605 ;
        RECT 175.285 47.995 175.455 48.165 ;
        RECT 175.285 42.555 175.455 42.725 ;
        RECT 175.285 37.115 175.455 37.285 ;
        RECT 175.285 31.675 175.455 31.845 ;
        RECT 175.285 26.235 175.455 26.405 ;
        RECT 175.285 20.795 175.455 20.965 ;
        RECT 175.285 15.355 175.455 15.525 ;
        RECT 175.285 9.915 175.455 10.085 ;
        RECT 175.745 58.875 175.915 59.045 ;
        RECT 175.745 53.435 175.915 53.605 ;
        RECT 175.745 47.995 175.915 48.165 ;
        RECT 175.745 42.555 175.915 42.725 ;
        RECT 175.745 37.115 175.915 37.285 ;
        RECT 175.745 31.675 175.915 31.845 ;
        RECT 175.745 26.235 175.915 26.405 ;
        RECT 175.745 20.795 175.915 20.965 ;
        RECT 175.745 15.355 175.915 15.525 ;
        RECT 175.745 9.915 175.915 10.085 ;
        RECT 176.205 58.875 176.375 59.045 ;
        RECT 176.205 53.435 176.375 53.605 ;
        RECT 176.205 47.995 176.375 48.165 ;
        RECT 176.205 42.555 176.375 42.725 ;
        RECT 176.205 37.115 176.375 37.285 ;
        RECT 176.205 31.675 176.375 31.845 ;
        RECT 176.205 26.235 176.375 26.405 ;
        RECT 176.205 20.795 176.375 20.965 ;
        RECT 176.205 15.355 176.375 15.525 ;
        RECT 176.205 9.915 176.375 10.085 ;
        RECT 176.665 58.875 176.835 59.045 ;
        RECT 176.665 53.435 176.835 53.605 ;
        RECT 176.665 47.995 176.835 48.165 ;
        RECT 176.665 42.555 176.835 42.725 ;
        RECT 176.665 37.115 176.835 37.285 ;
        RECT 176.665 31.675 176.835 31.845 ;
        RECT 176.665 26.235 176.835 26.405 ;
        RECT 176.665 20.795 176.835 20.965 ;
        RECT 176.665 15.355 176.835 15.525 ;
        RECT 176.665 9.915 176.835 10.085 ;
        RECT 177.125 58.875 177.295 59.045 ;
        RECT 177.125 53.435 177.295 53.605 ;
        RECT 177.125 47.995 177.295 48.165 ;
        RECT 177.125 42.555 177.295 42.725 ;
        RECT 177.125 37.115 177.295 37.285 ;
        RECT 177.125 31.675 177.295 31.845 ;
        RECT 177.125 26.235 177.295 26.405 ;
        RECT 177.125 20.795 177.295 20.965 ;
        RECT 177.125 15.355 177.295 15.525 ;
        RECT 177.125 9.915 177.295 10.085 ;
        RECT 177.585 58.875 177.755 59.045 ;
        RECT 177.585 53.435 177.755 53.605 ;
        RECT 177.585 47.995 177.755 48.165 ;
        RECT 177.585 42.555 177.755 42.725 ;
        RECT 177.585 37.115 177.755 37.285 ;
        RECT 177.585 31.675 177.755 31.845 ;
        RECT 177.585 26.235 177.755 26.405 ;
        RECT 177.585 20.795 177.755 20.965 ;
        RECT 177.585 15.355 177.755 15.525 ;
        RECT 177.585 9.915 177.755 10.085 ;
        RECT 178.045 58.875 178.215 59.045 ;
        RECT 178.045 53.435 178.215 53.605 ;
        RECT 178.045 47.995 178.215 48.165 ;
        RECT 178.045 42.555 178.215 42.725 ;
        RECT 178.045 37.115 178.215 37.285 ;
        RECT 178.045 31.675 178.215 31.845 ;
        RECT 178.045 26.235 178.215 26.405 ;
        RECT 178.045 20.795 178.215 20.965 ;
        RECT 178.045 15.355 178.215 15.525 ;
        RECT 178.045 9.915 178.215 10.085 ;
        RECT 178.505 58.875 178.675 59.045 ;
        RECT 178.505 53.435 178.675 53.605 ;
        RECT 178.505 47.995 178.675 48.165 ;
        RECT 178.505 42.555 178.675 42.725 ;
        RECT 178.505 37.115 178.675 37.285 ;
        RECT 178.505 31.675 178.675 31.845 ;
        RECT 178.505 26.235 178.675 26.405 ;
        RECT 178.505 20.795 178.675 20.965 ;
        RECT 178.505 15.355 178.675 15.525 ;
        RECT 178.505 9.915 178.675 10.085 ;
        RECT 178.965 58.875 179.135 59.045 ;
        RECT 178.965 53.435 179.135 53.605 ;
        RECT 178.965 47.995 179.135 48.165 ;
        RECT 178.965 42.555 179.135 42.725 ;
        RECT 178.965 37.115 179.135 37.285 ;
        RECT 178.965 31.675 179.135 31.845 ;
        RECT 178.965 26.235 179.135 26.405 ;
        RECT 178.965 20.795 179.135 20.965 ;
        RECT 178.965 15.355 179.135 15.525 ;
        RECT 178.965 9.915 179.135 10.085 ;
        RECT 179.425 58.875 179.595 59.045 ;
        RECT 179.425 53.435 179.595 53.605 ;
        RECT 179.425 47.995 179.595 48.165 ;
        RECT 179.425 42.555 179.595 42.725 ;
        RECT 179.425 37.115 179.595 37.285 ;
        RECT 179.425 31.675 179.595 31.845 ;
        RECT 179.425 26.235 179.595 26.405 ;
        RECT 179.425 20.795 179.595 20.965 ;
        RECT 179.425 15.355 179.595 15.525 ;
        RECT 179.425 9.915 179.595 10.085 ;
        RECT 179.885 58.875 180.055 59.045 ;
        RECT 179.885 53.435 180.055 53.605 ;
        RECT 179.885 47.995 180.055 48.165 ;
        RECT 179.885 42.555 180.055 42.725 ;
        RECT 179.885 37.115 180.055 37.285 ;
        RECT 179.885 31.675 180.055 31.845 ;
        RECT 179.885 26.235 180.055 26.405 ;
        RECT 179.885 20.795 180.055 20.965 ;
        RECT 179.885 15.355 180.055 15.525 ;
        RECT 179.885 9.915 180.055 10.085 ;
        RECT 180.345 58.875 180.515 59.045 ;
        RECT 180.345 53.435 180.515 53.605 ;
        RECT 180.345 47.995 180.515 48.165 ;
        RECT 180.345 42.555 180.515 42.725 ;
        RECT 180.345 37.115 180.515 37.285 ;
        RECT 180.345 31.675 180.515 31.845 ;
        RECT 180.345 26.235 180.515 26.405 ;
        RECT 180.345 20.795 180.515 20.965 ;
        RECT 180.345 15.355 180.515 15.525 ;
        RECT 180.345 9.915 180.515 10.085 ;
        RECT 180.805 58.875 180.975 59.045 ;
        RECT 180.805 53.435 180.975 53.605 ;
        RECT 180.805 47.995 180.975 48.165 ;
        RECT 180.805 42.555 180.975 42.725 ;
        RECT 180.805 37.115 180.975 37.285 ;
        RECT 180.805 31.675 180.975 31.845 ;
        RECT 180.805 26.235 180.975 26.405 ;
        RECT 180.805 20.795 180.975 20.965 ;
        RECT 180.805 15.355 180.975 15.525 ;
        RECT 180.805 9.915 180.975 10.085 ;
        RECT 181.265 58.875 181.435 59.045 ;
        RECT 181.265 53.435 181.435 53.605 ;
        RECT 181.265 47.995 181.435 48.165 ;
        RECT 181.265 42.555 181.435 42.725 ;
        RECT 181.265 37.115 181.435 37.285 ;
        RECT 181.265 31.675 181.435 31.845 ;
        RECT 181.265 26.235 181.435 26.405 ;
        RECT 181.265 20.795 181.435 20.965 ;
        RECT 181.265 15.355 181.435 15.525 ;
        RECT 181.265 9.915 181.435 10.085 ;
        RECT 181.725 58.875 181.895 59.045 ;
        RECT 181.725 53.435 181.895 53.605 ;
        RECT 181.725 47.995 181.895 48.165 ;
        RECT 181.725 42.555 181.895 42.725 ;
        RECT 181.725 37.115 181.895 37.285 ;
        RECT 181.725 31.675 181.895 31.845 ;
        RECT 181.725 26.235 181.895 26.405 ;
        RECT 181.725 20.795 181.895 20.965 ;
        RECT 181.725 15.355 181.895 15.525 ;
        RECT 181.725 9.915 181.895 10.085 ;
        RECT 182.185 58.875 182.355 59.045 ;
        RECT 182.185 53.435 182.355 53.605 ;
        RECT 182.185 47.995 182.355 48.165 ;
        RECT 182.185 42.555 182.355 42.725 ;
        RECT 182.185 37.115 182.355 37.285 ;
        RECT 182.185 31.675 182.355 31.845 ;
        RECT 182.185 26.235 182.355 26.405 ;
        RECT 182.185 20.795 182.355 20.965 ;
        RECT 182.185 15.355 182.355 15.525 ;
        RECT 182.185 9.915 182.355 10.085 ;
        RECT 182.645 58.875 182.815 59.045 ;
        RECT 182.645 53.435 182.815 53.605 ;
        RECT 182.645 47.995 182.815 48.165 ;
        RECT 182.645 42.555 182.815 42.725 ;
        RECT 182.645 37.115 182.815 37.285 ;
        RECT 182.645 31.675 182.815 31.845 ;
        RECT 182.645 26.235 182.815 26.405 ;
        RECT 182.645 20.795 182.815 20.965 ;
        RECT 182.645 15.355 182.815 15.525 ;
        RECT 182.645 9.915 182.815 10.085 ;
        RECT 183.105 58.875 183.275 59.045 ;
        RECT 183.105 53.435 183.275 53.605 ;
        RECT 183.105 47.995 183.275 48.165 ;
        RECT 183.105 42.555 183.275 42.725 ;
        RECT 183.105 37.115 183.275 37.285 ;
        RECT 183.105 31.675 183.275 31.845 ;
        RECT 183.105 26.235 183.275 26.405 ;
        RECT 183.105 20.795 183.275 20.965 ;
        RECT 183.105 15.355 183.275 15.525 ;
        RECT 183.105 9.915 183.275 10.085 ;
        RECT 183.565 58.875 183.735 59.045 ;
        RECT 183.565 53.435 183.735 53.605 ;
        RECT 183.565 47.995 183.735 48.165 ;
        RECT 183.565 42.555 183.735 42.725 ;
        RECT 183.565 37.115 183.735 37.285 ;
        RECT 183.565 31.675 183.735 31.845 ;
        RECT 183.565 26.235 183.735 26.405 ;
        RECT 183.565 20.795 183.735 20.965 ;
        RECT 183.565 15.355 183.735 15.525 ;
        RECT 183.565 9.915 183.735 10.085 ;
        RECT 184.025 58.875 184.195 59.045 ;
        RECT 184.025 53.435 184.195 53.605 ;
        RECT 184.025 47.995 184.195 48.165 ;
        RECT 184.025 42.555 184.195 42.725 ;
        RECT 184.025 37.115 184.195 37.285 ;
        RECT 184.025 31.675 184.195 31.845 ;
        RECT 184.025 26.235 184.195 26.405 ;
        RECT 184.025 20.795 184.195 20.965 ;
        RECT 184.025 15.355 184.195 15.525 ;
        RECT 184.025 9.915 184.195 10.085 ;
        RECT 184.485 58.875 184.655 59.045 ;
        RECT 184.485 53.435 184.655 53.605 ;
        RECT 184.485 47.995 184.655 48.165 ;
        RECT 184.485 42.555 184.655 42.725 ;
        RECT 184.485 37.115 184.655 37.285 ;
        RECT 184.485 31.675 184.655 31.845 ;
        RECT 184.485 26.235 184.655 26.405 ;
        RECT 184.485 20.795 184.655 20.965 ;
        RECT 184.485 15.355 184.655 15.525 ;
        RECT 184.485 9.915 184.655 10.085 ;
        RECT 184.945 58.875 185.115 59.045 ;
        RECT 184.945 53.435 185.115 53.605 ;
        RECT 184.945 47.995 185.115 48.165 ;
        RECT 184.945 42.555 185.115 42.725 ;
        RECT 184.945 37.115 185.115 37.285 ;
        RECT 184.945 31.675 185.115 31.845 ;
        RECT 184.945 26.235 185.115 26.405 ;
        RECT 184.945 20.795 185.115 20.965 ;
        RECT 184.945 15.355 185.115 15.525 ;
        RECT 184.945 9.915 185.115 10.085 ;
        RECT 185.405 58.875 185.575 59.045 ;
        RECT 185.405 53.435 185.575 53.605 ;
        RECT 185.405 47.995 185.575 48.165 ;
        RECT 185.405 42.555 185.575 42.725 ;
        RECT 185.405 37.115 185.575 37.285 ;
        RECT 185.405 31.675 185.575 31.845 ;
        RECT 185.405 26.235 185.575 26.405 ;
        RECT 185.405 20.795 185.575 20.965 ;
        RECT 185.405 15.355 185.575 15.525 ;
        RECT 185.405 9.915 185.575 10.085 ;
        RECT 185.865 58.875 186.035 59.045 ;
        RECT 185.865 53.435 186.035 53.605 ;
        RECT 185.865 47.995 186.035 48.165 ;
        RECT 185.865 42.555 186.035 42.725 ;
        RECT 185.865 37.115 186.035 37.285 ;
        RECT 185.865 31.675 186.035 31.845 ;
        RECT 185.865 26.235 186.035 26.405 ;
        RECT 185.865 20.795 186.035 20.965 ;
        RECT 185.865 15.355 186.035 15.525 ;
        RECT 185.865 9.915 186.035 10.085 ;
        RECT 186.325 58.875 186.495 59.045 ;
        RECT 186.325 53.435 186.495 53.605 ;
        RECT 186.325 47.995 186.495 48.165 ;
        RECT 186.325 42.555 186.495 42.725 ;
        RECT 186.325 37.115 186.495 37.285 ;
        RECT 186.325 31.675 186.495 31.845 ;
        RECT 186.325 26.235 186.495 26.405 ;
        RECT 186.325 20.795 186.495 20.965 ;
        RECT 186.325 15.355 186.495 15.525 ;
        RECT 186.325 9.915 186.495 10.085 ;
        RECT 186.785 58.875 186.955 59.045 ;
        RECT 186.785 53.435 186.955 53.605 ;
        RECT 186.785 47.995 186.955 48.165 ;
        RECT 186.785 42.555 186.955 42.725 ;
        RECT 186.785 37.115 186.955 37.285 ;
        RECT 186.785 31.675 186.955 31.845 ;
        RECT 186.785 26.235 186.955 26.405 ;
        RECT 186.785 20.795 186.955 20.965 ;
        RECT 186.785 15.355 186.955 15.525 ;
        RECT 186.785 9.915 186.955 10.085 ;
        RECT 187.245 58.875 187.415 59.045 ;
        RECT 187.245 53.435 187.415 53.605 ;
        RECT 187.245 47.995 187.415 48.165 ;
        RECT 187.245 42.555 187.415 42.725 ;
        RECT 187.245 37.115 187.415 37.285 ;
        RECT 187.245 31.675 187.415 31.845 ;
        RECT 187.245 26.235 187.415 26.405 ;
        RECT 187.245 20.795 187.415 20.965 ;
        RECT 187.245 15.355 187.415 15.525 ;
        RECT 187.245 9.915 187.415 10.085 ;
        RECT 187.705 58.875 187.875 59.045 ;
        RECT 187.705 53.435 187.875 53.605 ;
        RECT 187.705 47.995 187.875 48.165 ;
        RECT 187.705 42.555 187.875 42.725 ;
        RECT 187.705 37.115 187.875 37.285 ;
        RECT 187.705 31.675 187.875 31.845 ;
        RECT 187.705 26.235 187.875 26.405 ;
        RECT 187.705 20.795 187.875 20.965 ;
        RECT 187.705 15.355 187.875 15.525 ;
        RECT 187.705 9.915 187.875 10.085 ;
        RECT 188.165 58.875 188.335 59.045 ;
        RECT 188.165 53.435 188.335 53.605 ;
        RECT 188.165 47.995 188.335 48.165 ;
        RECT 188.165 42.555 188.335 42.725 ;
        RECT 188.165 37.115 188.335 37.285 ;
        RECT 188.165 31.675 188.335 31.845 ;
        RECT 188.165 26.235 188.335 26.405 ;
        RECT 188.165 20.795 188.335 20.965 ;
        RECT 188.165 15.355 188.335 15.525 ;
        RECT 188.165 9.915 188.335 10.085 ;
        RECT 188.625 58.875 188.795 59.045 ;
        RECT 188.625 53.435 188.795 53.605 ;
        RECT 188.625 47.995 188.795 48.165 ;
        RECT 188.625 42.555 188.795 42.725 ;
        RECT 188.625 37.115 188.795 37.285 ;
        RECT 188.625 31.675 188.795 31.845 ;
        RECT 188.625 26.235 188.795 26.405 ;
        RECT 188.625 20.795 188.795 20.965 ;
        RECT 188.625 15.355 188.795 15.525 ;
        RECT 188.625 9.915 188.795 10.085 ;
        RECT 189.085 58.875 189.255 59.045 ;
        RECT 189.085 53.435 189.255 53.605 ;
        RECT 189.085 47.995 189.255 48.165 ;
        RECT 189.085 42.555 189.255 42.725 ;
        RECT 189.085 37.115 189.255 37.285 ;
        RECT 189.085 31.675 189.255 31.845 ;
        RECT 189.085 26.235 189.255 26.405 ;
        RECT 189.085 20.795 189.255 20.965 ;
        RECT 189.085 15.355 189.255 15.525 ;
        RECT 189.085 9.915 189.255 10.085 ;
        RECT 189.545 58.875 189.715 59.045 ;
        RECT 189.545 53.435 189.715 53.605 ;
        RECT 189.545 47.995 189.715 48.165 ;
        RECT 189.545 42.555 189.715 42.725 ;
        RECT 189.545 37.115 189.715 37.285 ;
        RECT 189.545 31.675 189.715 31.845 ;
        RECT 189.545 26.235 189.715 26.405 ;
        RECT 189.545 20.795 189.715 20.965 ;
        RECT 189.545 15.355 189.715 15.525 ;
        RECT 189.545 9.915 189.715 10.085 ;
        RECT 102.145 58.875 102.315 59.045 ;
        RECT 102.145 53.435 102.315 53.605 ;
        RECT 102.145 47.995 102.315 48.165 ;
        RECT 102.145 42.555 102.315 42.725 ;
        RECT 102.145 37.115 102.315 37.285 ;
        RECT 102.145 31.675 102.315 31.845 ;
        RECT 102.145 26.235 102.315 26.405 ;
        RECT 102.145 20.795 102.315 20.965 ;
        RECT 102.145 15.355 102.315 15.525 ;
        RECT 102.145 9.915 102.315 10.085 ;
        RECT 102.605 58.875 102.775 59.045 ;
        RECT 102.605 53.435 102.775 53.605 ;
        RECT 102.605 47.995 102.775 48.165 ;
        RECT 102.605 42.555 102.775 42.725 ;
        RECT 102.605 37.115 102.775 37.285 ;
        RECT 102.605 31.675 102.775 31.845 ;
        RECT 102.605 26.235 102.775 26.405 ;
        RECT 102.605 20.795 102.775 20.965 ;
        RECT 102.605 15.355 102.775 15.525 ;
        RECT 102.605 9.915 102.775 10.085 ;
        RECT 103.065 58.875 103.235 59.045 ;
        RECT 103.065 53.435 103.235 53.605 ;
        RECT 103.065 47.995 103.235 48.165 ;
        RECT 103.065 42.555 103.235 42.725 ;
        RECT 103.065 37.115 103.235 37.285 ;
        RECT 103.065 31.675 103.235 31.845 ;
        RECT 103.065 26.235 103.235 26.405 ;
        RECT 103.065 20.795 103.235 20.965 ;
        RECT 103.065 15.355 103.235 15.525 ;
        RECT 103.065 9.915 103.235 10.085 ;
        RECT 103.525 58.875 103.695 59.045 ;
        RECT 103.525 53.435 103.695 53.605 ;
        RECT 103.525 47.995 103.695 48.165 ;
        RECT 103.525 42.555 103.695 42.725 ;
        RECT 103.525 37.115 103.695 37.285 ;
        RECT 103.525 31.675 103.695 31.845 ;
        RECT 103.525 26.235 103.695 26.405 ;
        RECT 103.525 20.795 103.695 20.965 ;
        RECT 103.525 15.355 103.695 15.525 ;
        RECT 103.525 9.915 103.695 10.085 ;
        RECT 103.985 58.875 104.155 59.045 ;
        RECT 103.985 53.435 104.155 53.605 ;
        RECT 103.985 47.995 104.155 48.165 ;
        RECT 103.985 42.555 104.155 42.725 ;
        RECT 103.985 37.115 104.155 37.285 ;
        RECT 103.985 31.675 104.155 31.845 ;
        RECT 103.985 26.235 104.155 26.405 ;
        RECT 103.985 20.795 104.155 20.965 ;
        RECT 103.985 15.355 104.155 15.525 ;
        RECT 103.985 9.915 104.155 10.085 ;
        RECT 104.445 58.875 104.615 59.045 ;
        RECT 104.445 53.435 104.615 53.605 ;
        RECT 104.445 47.995 104.615 48.165 ;
        RECT 104.445 42.555 104.615 42.725 ;
        RECT 104.445 37.115 104.615 37.285 ;
        RECT 104.445 31.675 104.615 31.845 ;
        RECT 104.445 26.235 104.615 26.405 ;
        RECT 104.445 20.795 104.615 20.965 ;
        RECT 104.445 15.355 104.615 15.525 ;
        RECT 104.445 9.915 104.615 10.085 ;
        RECT 104.905 58.875 105.075 59.045 ;
        RECT 104.905 53.435 105.075 53.605 ;
        RECT 104.905 47.995 105.075 48.165 ;
        RECT 104.905 42.555 105.075 42.725 ;
        RECT 104.905 37.115 105.075 37.285 ;
        RECT 104.905 31.675 105.075 31.845 ;
        RECT 104.905 26.235 105.075 26.405 ;
        RECT 104.905 20.795 105.075 20.965 ;
        RECT 104.905 15.355 105.075 15.525 ;
        RECT 104.905 9.915 105.075 10.085 ;
        RECT 105.365 58.875 105.535 59.045 ;
        RECT 105.365 53.435 105.535 53.605 ;
        RECT 105.365 47.995 105.535 48.165 ;
        RECT 105.365 42.555 105.535 42.725 ;
        RECT 105.365 37.115 105.535 37.285 ;
        RECT 105.365 31.675 105.535 31.845 ;
        RECT 105.365 26.235 105.535 26.405 ;
        RECT 105.365 20.795 105.535 20.965 ;
        RECT 105.365 15.355 105.535 15.525 ;
        RECT 105.365 9.915 105.535 10.085 ;
        RECT 105.825 58.875 105.995 59.045 ;
        RECT 105.825 53.435 105.995 53.605 ;
        RECT 105.825 47.995 105.995 48.165 ;
        RECT 105.825 42.555 105.995 42.725 ;
        RECT 105.825 37.115 105.995 37.285 ;
        RECT 105.825 31.675 105.995 31.845 ;
        RECT 105.825 26.235 105.995 26.405 ;
        RECT 105.825 20.795 105.995 20.965 ;
        RECT 105.825 15.355 105.995 15.525 ;
        RECT 105.825 9.915 105.995 10.085 ;
        RECT 106.285 58.875 106.455 59.045 ;
        RECT 106.285 53.435 106.455 53.605 ;
        RECT 106.285 47.995 106.455 48.165 ;
        RECT 106.285 42.555 106.455 42.725 ;
        RECT 106.285 37.115 106.455 37.285 ;
        RECT 106.285 31.675 106.455 31.845 ;
        RECT 106.285 26.235 106.455 26.405 ;
        RECT 106.285 20.795 106.455 20.965 ;
        RECT 106.285 15.355 106.455 15.525 ;
        RECT 106.285 9.915 106.455 10.085 ;
        RECT 106.745 58.875 106.915 59.045 ;
        RECT 106.745 53.435 106.915 53.605 ;
        RECT 106.745 47.995 106.915 48.165 ;
        RECT 106.745 42.555 106.915 42.725 ;
        RECT 106.745 37.115 106.915 37.285 ;
        RECT 106.745 31.675 106.915 31.845 ;
        RECT 106.745 26.235 106.915 26.405 ;
        RECT 106.745 20.795 106.915 20.965 ;
        RECT 106.745 15.355 106.915 15.525 ;
        RECT 106.745 9.915 106.915 10.085 ;
        RECT 107.205 58.875 107.375 59.045 ;
        RECT 107.205 53.435 107.375 53.605 ;
        RECT 107.205 47.995 107.375 48.165 ;
        RECT 107.205 42.555 107.375 42.725 ;
        RECT 107.205 37.115 107.375 37.285 ;
        RECT 107.205 31.675 107.375 31.845 ;
        RECT 107.205 26.235 107.375 26.405 ;
        RECT 107.205 20.795 107.375 20.965 ;
        RECT 107.205 15.355 107.375 15.525 ;
        RECT 107.205 9.915 107.375 10.085 ;
        RECT 107.665 58.875 107.835 59.045 ;
        RECT 107.665 53.435 107.835 53.605 ;
        RECT 107.665 47.995 107.835 48.165 ;
        RECT 107.665 42.555 107.835 42.725 ;
        RECT 107.665 37.115 107.835 37.285 ;
        RECT 107.665 31.675 107.835 31.845 ;
        RECT 107.665 26.235 107.835 26.405 ;
        RECT 107.665 20.795 107.835 20.965 ;
        RECT 107.665 15.355 107.835 15.525 ;
        RECT 107.665 9.915 107.835 10.085 ;
        RECT 108.125 58.875 108.295 59.045 ;
        RECT 108.125 53.435 108.295 53.605 ;
        RECT 108.125 47.995 108.295 48.165 ;
        RECT 108.125 42.555 108.295 42.725 ;
        RECT 108.125 37.115 108.295 37.285 ;
        RECT 108.125 31.675 108.295 31.845 ;
        RECT 108.125 26.235 108.295 26.405 ;
        RECT 108.125 20.795 108.295 20.965 ;
        RECT 108.125 15.355 108.295 15.525 ;
        RECT 108.125 9.915 108.295 10.085 ;
        RECT 108.585 58.875 108.755 59.045 ;
        RECT 108.585 53.435 108.755 53.605 ;
        RECT 108.585 47.995 108.755 48.165 ;
        RECT 108.585 42.555 108.755 42.725 ;
        RECT 108.585 37.115 108.755 37.285 ;
        RECT 108.585 31.675 108.755 31.845 ;
        RECT 108.585 26.235 108.755 26.405 ;
        RECT 108.585 20.795 108.755 20.965 ;
        RECT 108.585 15.355 108.755 15.525 ;
        RECT 108.585 9.915 108.755 10.085 ;
        RECT 109.045 58.875 109.215 59.045 ;
        RECT 109.045 53.435 109.215 53.605 ;
        RECT 109.045 47.995 109.215 48.165 ;
        RECT 109.045 42.555 109.215 42.725 ;
        RECT 109.045 37.115 109.215 37.285 ;
        RECT 109.045 31.675 109.215 31.845 ;
        RECT 109.045 26.235 109.215 26.405 ;
        RECT 109.045 20.795 109.215 20.965 ;
        RECT 109.045 15.355 109.215 15.525 ;
        RECT 109.045 9.915 109.215 10.085 ;
        RECT 109.505 58.875 109.675 59.045 ;
        RECT 109.505 53.435 109.675 53.605 ;
        RECT 109.505 47.995 109.675 48.165 ;
        RECT 109.505 42.555 109.675 42.725 ;
        RECT 109.505 37.115 109.675 37.285 ;
        RECT 109.505 31.675 109.675 31.845 ;
        RECT 109.505 26.235 109.675 26.405 ;
        RECT 109.505 20.795 109.675 20.965 ;
        RECT 109.505 15.355 109.675 15.525 ;
        RECT 109.505 9.915 109.675 10.085 ;
        RECT 109.965 58.875 110.135 59.045 ;
        RECT 109.965 53.435 110.135 53.605 ;
        RECT 109.965 47.995 110.135 48.165 ;
        RECT 109.965 42.555 110.135 42.725 ;
        RECT 109.965 37.115 110.135 37.285 ;
        RECT 109.965 31.675 110.135 31.845 ;
        RECT 109.965 26.235 110.135 26.405 ;
        RECT 109.965 20.795 110.135 20.965 ;
        RECT 109.965 15.355 110.135 15.525 ;
        RECT 109.965 9.915 110.135 10.085 ;
        RECT 110.425 58.875 110.595 59.045 ;
        RECT 110.425 53.435 110.595 53.605 ;
        RECT 110.425 47.995 110.595 48.165 ;
        RECT 110.425 42.555 110.595 42.725 ;
        RECT 110.425 37.115 110.595 37.285 ;
        RECT 110.425 31.675 110.595 31.845 ;
        RECT 110.425 26.235 110.595 26.405 ;
        RECT 110.425 20.795 110.595 20.965 ;
        RECT 110.425 15.355 110.595 15.525 ;
        RECT 110.425 9.915 110.595 10.085 ;
        RECT 110.885 58.875 111.055 59.045 ;
        RECT 110.885 53.435 111.055 53.605 ;
        RECT 110.885 47.995 111.055 48.165 ;
        RECT 110.885 42.555 111.055 42.725 ;
        RECT 110.885 37.115 111.055 37.285 ;
        RECT 110.885 31.675 111.055 31.845 ;
        RECT 110.885 26.235 111.055 26.405 ;
        RECT 110.885 20.795 111.055 20.965 ;
        RECT 110.885 15.355 111.055 15.525 ;
        RECT 110.885 9.915 111.055 10.085 ;
        RECT 111.345 58.875 111.515 59.045 ;
        RECT 111.345 53.435 111.515 53.605 ;
        RECT 111.345 47.995 111.515 48.165 ;
        RECT 111.345 42.555 111.515 42.725 ;
        RECT 111.345 37.115 111.515 37.285 ;
        RECT 111.345 31.675 111.515 31.845 ;
        RECT 111.345 26.235 111.515 26.405 ;
        RECT 111.345 20.795 111.515 20.965 ;
        RECT 111.345 15.355 111.515 15.525 ;
        RECT 111.345 9.915 111.515 10.085 ;
        RECT 111.805 58.875 111.975 59.045 ;
        RECT 111.805 53.435 111.975 53.605 ;
        RECT 111.805 47.995 111.975 48.165 ;
        RECT 111.805 42.555 111.975 42.725 ;
        RECT 111.805 37.115 111.975 37.285 ;
        RECT 111.805 31.675 111.975 31.845 ;
        RECT 111.805 26.235 111.975 26.405 ;
        RECT 111.805 20.795 111.975 20.965 ;
        RECT 111.805 15.355 111.975 15.525 ;
        RECT 111.805 9.915 111.975 10.085 ;
        RECT 112.265 58.875 112.435 59.045 ;
        RECT 112.265 53.435 112.435 53.605 ;
        RECT 112.265 47.995 112.435 48.165 ;
        RECT 112.265 42.555 112.435 42.725 ;
        RECT 112.265 37.115 112.435 37.285 ;
        RECT 112.265 31.675 112.435 31.845 ;
        RECT 112.265 26.235 112.435 26.405 ;
        RECT 112.265 20.795 112.435 20.965 ;
        RECT 112.265 15.355 112.435 15.525 ;
        RECT 112.265 9.915 112.435 10.085 ;
        RECT 112.725 58.875 112.895 59.045 ;
        RECT 112.725 53.435 112.895 53.605 ;
        RECT 112.725 47.995 112.895 48.165 ;
        RECT 112.725 42.555 112.895 42.725 ;
        RECT 112.725 37.115 112.895 37.285 ;
        RECT 112.725 31.675 112.895 31.845 ;
        RECT 112.725 26.235 112.895 26.405 ;
        RECT 112.725 20.795 112.895 20.965 ;
        RECT 112.725 15.355 112.895 15.525 ;
        RECT 112.725 9.915 112.895 10.085 ;
        RECT 113.185 58.875 113.355 59.045 ;
        RECT 113.185 53.435 113.355 53.605 ;
        RECT 113.185 47.995 113.355 48.165 ;
        RECT 113.185 42.555 113.355 42.725 ;
        RECT 113.185 37.115 113.355 37.285 ;
        RECT 113.185 31.675 113.355 31.845 ;
        RECT 113.185 26.235 113.355 26.405 ;
        RECT 113.185 20.795 113.355 20.965 ;
        RECT 113.185 15.355 113.355 15.525 ;
        RECT 113.185 9.915 113.355 10.085 ;
        RECT 113.645 58.875 113.815 59.045 ;
        RECT 113.645 53.435 113.815 53.605 ;
        RECT 113.645 47.995 113.815 48.165 ;
        RECT 113.645 42.555 113.815 42.725 ;
        RECT 113.645 37.115 113.815 37.285 ;
        RECT 113.645 31.675 113.815 31.845 ;
        RECT 113.645 26.235 113.815 26.405 ;
        RECT 113.645 20.795 113.815 20.965 ;
        RECT 113.645 15.355 113.815 15.525 ;
        RECT 113.645 9.915 113.815 10.085 ;
        RECT 114.105 58.875 114.275 59.045 ;
        RECT 114.105 53.435 114.275 53.605 ;
        RECT 114.105 47.995 114.275 48.165 ;
        RECT 114.105 42.555 114.275 42.725 ;
        RECT 114.105 37.115 114.275 37.285 ;
        RECT 114.105 31.675 114.275 31.845 ;
        RECT 114.105 26.235 114.275 26.405 ;
        RECT 114.105 20.795 114.275 20.965 ;
        RECT 114.105 15.355 114.275 15.525 ;
        RECT 114.105 9.915 114.275 10.085 ;
        RECT 114.565 58.875 114.735 59.045 ;
        RECT 114.565 53.435 114.735 53.605 ;
        RECT 114.565 47.995 114.735 48.165 ;
        RECT 114.565 42.555 114.735 42.725 ;
        RECT 114.565 37.115 114.735 37.285 ;
        RECT 114.565 31.675 114.735 31.845 ;
        RECT 114.565 26.235 114.735 26.405 ;
        RECT 114.565 20.795 114.735 20.965 ;
        RECT 114.565 15.355 114.735 15.525 ;
        RECT 114.565 9.915 114.735 10.085 ;
        RECT 115.025 58.875 115.195 59.045 ;
        RECT 115.025 53.435 115.195 53.605 ;
        RECT 115.025 47.995 115.195 48.165 ;
        RECT 115.025 42.555 115.195 42.725 ;
        RECT 115.025 37.115 115.195 37.285 ;
        RECT 115.025 31.675 115.195 31.845 ;
        RECT 115.025 26.235 115.195 26.405 ;
        RECT 115.025 20.795 115.195 20.965 ;
        RECT 115.025 15.355 115.195 15.525 ;
        RECT 115.025 9.915 115.195 10.085 ;
        RECT 115.485 58.875 115.655 59.045 ;
        RECT 115.485 53.435 115.655 53.605 ;
        RECT 115.485 47.995 115.655 48.165 ;
        RECT 115.485 42.555 115.655 42.725 ;
        RECT 115.485 37.115 115.655 37.285 ;
        RECT 115.485 31.675 115.655 31.845 ;
        RECT 115.485 26.235 115.655 26.405 ;
        RECT 115.485 20.795 115.655 20.965 ;
        RECT 115.485 15.355 115.655 15.525 ;
        RECT 115.485 9.915 115.655 10.085 ;
        RECT 115.945 58.875 116.115 59.045 ;
        RECT 115.945 53.435 116.115 53.605 ;
        RECT 115.945 47.995 116.115 48.165 ;
        RECT 115.945 42.555 116.115 42.725 ;
        RECT 115.945 37.115 116.115 37.285 ;
        RECT 115.945 31.675 116.115 31.845 ;
        RECT 115.945 26.235 116.115 26.405 ;
        RECT 115.945 20.795 116.115 20.965 ;
        RECT 115.945 15.355 116.115 15.525 ;
        RECT 115.945 9.915 116.115 10.085 ;
        RECT 116.405 58.875 116.575 59.045 ;
        RECT 116.405 53.435 116.575 53.605 ;
        RECT 116.405 47.995 116.575 48.165 ;
        RECT 116.405 42.555 116.575 42.725 ;
        RECT 116.405 37.115 116.575 37.285 ;
        RECT 116.405 31.675 116.575 31.845 ;
        RECT 116.405 26.235 116.575 26.405 ;
        RECT 116.405 20.795 116.575 20.965 ;
        RECT 116.405 15.355 116.575 15.525 ;
        RECT 116.405 9.915 116.575 10.085 ;
        RECT 116.865 58.875 117.035 59.045 ;
        RECT 116.865 53.435 117.035 53.605 ;
        RECT 116.865 47.995 117.035 48.165 ;
        RECT 116.865 42.555 117.035 42.725 ;
        RECT 116.865 37.115 117.035 37.285 ;
        RECT 116.865 31.675 117.035 31.845 ;
        RECT 116.865 26.235 117.035 26.405 ;
        RECT 116.865 20.795 117.035 20.965 ;
        RECT 116.865 15.355 117.035 15.525 ;
        RECT 116.865 9.915 117.035 10.085 ;
        RECT 117.325 58.875 117.495 59.045 ;
        RECT 117.325 53.435 117.495 53.605 ;
        RECT 117.325 47.995 117.495 48.165 ;
        RECT 117.325 42.555 117.495 42.725 ;
        RECT 117.325 37.115 117.495 37.285 ;
        RECT 117.325 31.675 117.495 31.845 ;
        RECT 117.325 26.235 117.495 26.405 ;
        RECT 117.325 20.795 117.495 20.965 ;
        RECT 117.325 15.355 117.495 15.525 ;
        RECT 117.325 9.915 117.495 10.085 ;
        RECT 117.785 58.875 117.955 59.045 ;
        RECT 117.785 53.435 117.955 53.605 ;
        RECT 117.785 47.995 117.955 48.165 ;
        RECT 117.785 42.555 117.955 42.725 ;
        RECT 117.785 37.115 117.955 37.285 ;
        RECT 117.785 31.675 117.955 31.845 ;
        RECT 117.785 26.235 117.955 26.405 ;
        RECT 117.785 20.795 117.955 20.965 ;
        RECT 117.785 15.355 117.955 15.525 ;
        RECT 117.785 9.915 117.955 10.085 ;
        RECT 118.245 58.875 118.415 59.045 ;
        RECT 118.245 53.435 118.415 53.605 ;
        RECT 118.245 47.995 118.415 48.165 ;
        RECT 118.245 42.555 118.415 42.725 ;
        RECT 118.245 37.115 118.415 37.285 ;
        RECT 118.245 31.675 118.415 31.845 ;
        RECT 118.245 26.235 118.415 26.405 ;
        RECT 118.245 20.795 118.415 20.965 ;
        RECT 118.245 15.355 118.415 15.525 ;
        RECT 118.245 9.915 118.415 10.085 ;
        RECT 118.705 58.875 118.875 59.045 ;
        RECT 118.705 53.435 118.875 53.605 ;
        RECT 118.705 47.995 118.875 48.165 ;
        RECT 118.705 42.555 118.875 42.725 ;
        RECT 118.705 37.115 118.875 37.285 ;
        RECT 118.705 31.675 118.875 31.845 ;
        RECT 118.705 26.235 118.875 26.405 ;
        RECT 118.705 20.795 118.875 20.965 ;
        RECT 118.705 15.355 118.875 15.525 ;
        RECT 118.705 9.915 118.875 10.085 ;
        RECT 119.165 58.875 119.335 59.045 ;
        RECT 119.165 53.435 119.335 53.605 ;
        RECT 119.165 47.995 119.335 48.165 ;
        RECT 119.165 42.555 119.335 42.725 ;
        RECT 119.165 37.115 119.335 37.285 ;
        RECT 119.165 31.675 119.335 31.845 ;
        RECT 119.165 26.235 119.335 26.405 ;
        RECT 119.165 20.795 119.335 20.965 ;
        RECT 119.165 15.355 119.335 15.525 ;
        RECT 119.165 9.915 119.335 10.085 ;
        RECT 119.625 58.875 119.795 59.045 ;
        RECT 119.625 53.435 119.795 53.605 ;
        RECT 119.625 47.995 119.795 48.165 ;
        RECT 119.625 42.555 119.795 42.725 ;
        RECT 119.625 37.115 119.795 37.285 ;
        RECT 119.625 31.675 119.795 31.845 ;
        RECT 119.625 26.235 119.795 26.405 ;
        RECT 119.625 20.795 119.795 20.965 ;
        RECT 119.625 15.355 119.795 15.525 ;
        RECT 119.625 9.915 119.795 10.085 ;
        RECT 120.085 58.875 120.255 59.045 ;
        RECT 120.085 53.435 120.255 53.605 ;
        RECT 120.085 47.995 120.255 48.165 ;
        RECT 120.085 42.555 120.255 42.725 ;
        RECT 120.085 37.115 120.255 37.285 ;
        RECT 120.085 31.675 120.255 31.845 ;
        RECT 120.085 26.235 120.255 26.405 ;
        RECT 120.085 20.795 120.255 20.965 ;
        RECT 120.085 15.355 120.255 15.525 ;
        RECT 120.085 9.915 120.255 10.085 ;
        RECT 120.545 58.875 120.715 59.045 ;
        RECT 120.545 53.435 120.715 53.605 ;
        RECT 120.545 47.995 120.715 48.165 ;
        RECT 120.545 42.555 120.715 42.725 ;
        RECT 120.545 37.115 120.715 37.285 ;
        RECT 120.545 31.675 120.715 31.845 ;
        RECT 120.545 26.235 120.715 26.405 ;
        RECT 120.545 20.795 120.715 20.965 ;
        RECT 120.545 15.355 120.715 15.525 ;
        RECT 120.545 9.915 120.715 10.085 ;
        RECT 121.005 58.875 121.175 59.045 ;
        RECT 121.005 53.435 121.175 53.605 ;
        RECT 121.005 47.995 121.175 48.165 ;
        RECT 121.005 42.555 121.175 42.725 ;
        RECT 121.005 37.115 121.175 37.285 ;
        RECT 121.005 31.675 121.175 31.845 ;
        RECT 121.005 26.235 121.175 26.405 ;
        RECT 121.005 20.795 121.175 20.965 ;
        RECT 121.005 15.355 121.175 15.525 ;
        RECT 121.005 9.915 121.175 10.085 ;
        RECT 121.465 58.875 121.635 59.045 ;
        RECT 121.465 53.435 121.635 53.605 ;
        RECT 121.465 47.995 121.635 48.165 ;
        RECT 121.465 42.555 121.635 42.725 ;
        RECT 121.465 37.115 121.635 37.285 ;
        RECT 121.465 31.675 121.635 31.845 ;
        RECT 121.465 26.235 121.635 26.405 ;
        RECT 121.465 20.795 121.635 20.965 ;
        RECT 121.465 15.355 121.635 15.525 ;
        RECT 121.465 9.915 121.635 10.085 ;
        RECT 121.925 58.875 122.095 59.045 ;
        RECT 121.925 53.435 122.095 53.605 ;
        RECT 121.925 47.995 122.095 48.165 ;
        RECT 121.925 42.555 122.095 42.725 ;
        RECT 121.925 37.115 122.095 37.285 ;
        RECT 121.925 31.675 122.095 31.845 ;
        RECT 121.925 26.235 122.095 26.405 ;
        RECT 121.925 20.795 122.095 20.965 ;
        RECT 121.925 15.355 122.095 15.525 ;
        RECT 121.925 9.915 122.095 10.085 ;
        RECT 122.385 58.875 122.555 59.045 ;
        RECT 122.385 53.435 122.555 53.605 ;
        RECT 122.385 47.995 122.555 48.165 ;
        RECT 122.385 42.555 122.555 42.725 ;
        RECT 122.385 37.115 122.555 37.285 ;
        RECT 122.385 31.675 122.555 31.845 ;
        RECT 122.385 26.235 122.555 26.405 ;
        RECT 122.385 20.795 122.555 20.965 ;
        RECT 122.385 15.355 122.555 15.525 ;
        RECT 122.385 9.915 122.555 10.085 ;
        RECT 122.845 58.875 123.015 59.045 ;
        RECT 122.845 53.435 123.015 53.605 ;
        RECT 122.845 47.995 123.015 48.165 ;
        RECT 122.845 42.555 123.015 42.725 ;
        RECT 122.845 37.115 123.015 37.285 ;
        RECT 122.845 31.675 123.015 31.845 ;
        RECT 122.845 26.235 123.015 26.405 ;
        RECT 122.845 20.795 123.015 20.965 ;
        RECT 122.845 15.355 123.015 15.525 ;
        RECT 122.845 9.915 123.015 10.085 ;
        RECT 123.305 58.875 123.475 59.045 ;
        RECT 123.305 53.435 123.475 53.605 ;
        RECT 123.305 47.995 123.475 48.165 ;
        RECT 123.305 42.555 123.475 42.725 ;
        RECT 123.305 37.115 123.475 37.285 ;
        RECT 123.305 31.675 123.475 31.845 ;
        RECT 123.305 26.235 123.475 26.405 ;
        RECT 123.305 20.795 123.475 20.965 ;
        RECT 123.305 15.355 123.475 15.525 ;
        RECT 123.305 9.915 123.475 10.085 ;
        RECT 123.765 58.875 123.935 59.045 ;
        RECT 123.765 53.435 123.935 53.605 ;
        RECT 123.765 47.995 123.935 48.165 ;
        RECT 123.765 42.555 123.935 42.725 ;
        RECT 123.765 37.115 123.935 37.285 ;
        RECT 123.765 31.675 123.935 31.845 ;
        RECT 123.765 26.235 123.935 26.405 ;
        RECT 123.765 20.795 123.935 20.965 ;
        RECT 123.765 15.355 123.935 15.525 ;
        RECT 123.765 9.915 123.935 10.085 ;
        RECT 124.225 58.875 124.395 59.045 ;
        RECT 124.225 53.435 124.395 53.605 ;
        RECT 124.225 47.995 124.395 48.165 ;
        RECT 124.225 42.555 124.395 42.725 ;
        RECT 124.225 37.115 124.395 37.285 ;
        RECT 124.225 31.675 124.395 31.845 ;
        RECT 124.225 26.235 124.395 26.405 ;
        RECT 124.225 20.795 124.395 20.965 ;
        RECT 124.225 15.355 124.395 15.525 ;
        RECT 124.225 9.915 124.395 10.085 ;
        RECT 124.685 58.875 124.855 59.045 ;
        RECT 124.685 53.435 124.855 53.605 ;
        RECT 124.685 47.995 124.855 48.165 ;
        RECT 124.685 42.555 124.855 42.725 ;
        RECT 124.685 37.115 124.855 37.285 ;
        RECT 124.685 31.675 124.855 31.845 ;
        RECT 124.685 26.235 124.855 26.405 ;
        RECT 124.685 20.795 124.855 20.965 ;
        RECT 124.685 15.355 124.855 15.525 ;
        RECT 124.685 9.915 124.855 10.085 ;
        RECT 125.145 58.875 125.315 59.045 ;
        RECT 125.145 53.435 125.315 53.605 ;
        RECT 125.145 47.995 125.315 48.165 ;
        RECT 125.145 42.555 125.315 42.725 ;
        RECT 125.145 37.115 125.315 37.285 ;
        RECT 125.145 31.675 125.315 31.845 ;
        RECT 125.145 26.235 125.315 26.405 ;
        RECT 125.145 20.795 125.315 20.965 ;
        RECT 125.145 15.355 125.315 15.525 ;
        RECT 125.145 9.915 125.315 10.085 ;
        RECT 125.605 58.875 125.775 59.045 ;
        RECT 125.605 53.435 125.775 53.605 ;
        RECT 125.605 47.995 125.775 48.165 ;
        RECT 125.605 42.555 125.775 42.725 ;
        RECT 125.605 37.115 125.775 37.285 ;
        RECT 125.605 31.675 125.775 31.845 ;
        RECT 125.605 26.235 125.775 26.405 ;
        RECT 125.605 20.795 125.775 20.965 ;
        RECT 125.605 15.355 125.775 15.525 ;
        RECT 125.605 9.915 125.775 10.085 ;
        RECT 126.065 58.875 126.235 59.045 ;
        RECT 126.065 53.435 126.235 53.605 ;
        RECT 126.065 47.995 126.235 48.165 ;
        RECT 126.065 42.555 126.235 42.725 ;
        RECT 126.065 37.115 126.235 37.285 ;
        RECT 126.065 31.675 126.235 31.845 ;
        RECT 126.065 26.235 126.235 26.405 ;
        RECT 126.065 20.795 126.235 20.965 ;
        RECT 126.065 15.355 126.235 15.525 ;
        RECT 126.065 9.915 126.235 10.085 ;
        RECT 126.525 58.875 126.695 59.045 ;
        RECT 126.525 53.435 126.695 53.605 ;
        RECT 126.525 47.995 126.695 48.165 ;
        RECT 126.525 42.555 126.695 42.725 ;
        RECT 126.525 37.115 126.695 37.285 ;
        RECT 126.525 31.675 126.695 31.845 ;
        RECT 126.525 26.235 126.695 26.405 ;
        RECT 126.525 20.795 126.695 20.965 ;
        RECT 126.525 15.355 126.695 15.525 ;
        RECT 126.525 9.915 126.695 10.085 ;
        RECT 126.985 58.875 127.155 59.045 ;
        RECT 126.985 53.435 127.155 53.605 ;
        RECT 126.985 47.995 127.155 48.165 ;
        RECT 126.985 42.555 127.155 42.725 ;
        RECT 126.985 37.115 127.155 37.285 ;
        RECT 126.985 31.675 127.155 31.845 ;
        RECT 126.985 26.235 127.155 26.405 ;
        RECT 126.985 20.795 127.155 20.965 ;
        RECT 126.985 15.355 127.155 15.525 ;
        RECT 126.985 9.915 127.155 10.085 ;
        RECT 127.445 58.875 127.615 59.045 ;
        RECT 127.445 53.435 127.615 53.605 ;
        RECT 127.445 47.995 127.615 48.165 ;
        RECT 127.445 42.555 127.615 42.725 ;
        RECT 127.445 37.115 127.615 37.285 ;
        RECT 127.445 31.675 127.615 31.845 ;
        RECT 127.445 26.235 127.615 26.405 ;
        RECT 127.445 20.795 127.615 20.965 ;
        RECT 127.445 15.355 127.615 15.525 ;
        RECT 127.445 9.915 127.615 10.085 ;
        RECT 127.905 58.875 128.075 59.045 ;
        RECT 127.905 53.435 128.075 53.605 ;
        RECT 127.905 47.995 128.075 48.165 ;
        RECT 127.905 42.555 128.075 42.725 ;
        RECT 127.905 37.115 128.075 37.285 ;
        RECT 127.905 31.675 128.075 31.845 ;
        RECT 127.905 26.235 128.075 26.405 ;
        RECT 127.905 20.795 128.075 20.965 ;
        RECT 127.905 15.355 128.075 15.525 ;
        RECT 127.905 9.915 128.075 10.085 ;
        RECT 128.365 58.875 128.535 59.045 ;
        RECT 128.365 53.435 128.535 53.605 ;
        RECT 128.365 47.995 128.535 48.165 ;
        RECT 128.365 42.555 128.535 42.725 ;
        RECT 128.365 37.115 128.535 37.285 ;
        RECT 128.365 31.675 128.535 31.845 ;
        RECT 128.365 26.235 128.535 26.405 ;
        RECT 128.365 20.795 128.535 20.965 ;
        RECT 128.365 15.355 128.535 15.525 ;
        RECT 128.365 9.915 128.535 10.085 ;
        RECT 128.825 58.875 128.995 59.045 ;
        RECT 128.825 53.435 128.995 53.605 ;
        RECT 128.825 47.995 128.995 48.165 ;
        RECT 128.825 42.555 128.995 42.725 ;
        RECT 128.825 37.115 128.995 37.285 ;
        RECT 128.825 31.675 128.995 31.845 ;
        RECT 128.825 26.235 128.995 26.405 ;
        RECT 128.825 20.795 128.995 20.965 ;
        RECT 128.825 15.355 128.995 15.525 ;
        RECT 128.825 9.915 128.995 10.085 ;
        RECT 129.285 58.875 129.455 59.045 ;
        RECT 129.285 53.435 129.455 53.605 ;
        RECT 129.285 47.995 129.455 48.165 ;
        RECT 129.285 42.555 129.455 42.725 ;
        RECT 129.285 37.115 129.455 37.285 ;
        RECT 129.285 31.675 129.455 31.845 ;
        RECT 129.285 26.235 129.455 26.405 ;
        RECT 129.285 20.795 129.455 20.965 ;
        RECT 129.285 15.355 129.455 15.525 ;
        RECT 129.285 9.915 129.455 10.085 ;
        RECT 129.745 58.875 129.915 59.045 ;
        RECT 129.745 53.435 129.915 53.605 ;
        RECT 129.745 47.995 129.915 48.165 ;
        RECT 129.745 42.555 129.915 42.725 ;
        RECT 129.745 37.115 129.915 37.285 ;
        RECT 129.745 31.675 129.915 31.845 ;
        RECT 129.745 26.235 129.915 26.405 ;
        RECT 129.745 20.795 129.915 20.965 ;
        RECT 129.745 15.355 129.915 15.525 ;
        RECT 129.745 9.915 129.915 10.085 ;
        RECT 130.205 58.875 130.375 59.045 ;
        RECT 130.205 53.435 130.375 53.605 ;
        RECT 130.205 47.995 130.375 48.165 ;
        RECT 130.205 42.555 130.375 42.725 ;
        RECT 130.205 37.115 130.375 37.285 ;
        RECT 130.205 31.675 130.375 31.845 ;
        RECT 130.205 26.235 130.375 26.405 ;
        RECT 130.205 20.795 130.375 20.965 ;
        RECT 130.205 15.355 130.375 15.525 ;
        RECT 130.205 9.915 130.375 10.085 ;
        RECT 130.665 58.875 130.835 59.045 ;
        RECT 130.665 53.435 130.835 53.605 ;
        RECT 130.665 47.995 130.835 48.165 ;
        RECT 130.665 42.555 130.835 42.725 ;
        RECT 130.665 37.115 130.835 37.285 ;
        RECT 130.665 31.675 130.835 31.845 ;
        RECT 130.665 26.235 130.835 26.405 ;
        RECT 130.665 20.795 130.835 20.965 ;
        RECT 130.665 15.355 130.835 15.525 ;
        RECT 130.665 9.915 130.835 10.085 ;
        RECT 131.125 58.875 131.295 59.045 ;
        RECT 131.125 53.435 131.295 53.605 ;
        RECT 131.125 47.995 131.295 48.165 ;
        RECT 131.125 42.555 131.295 42.725 ;
        RECT 131.125 37.115 131.295 37.285 ;
        RECT 131.125 31.675 131.295 31.845 ;
        RECT 131.125 26.235 131.295 26.405 ;
        RECT 131.125 20.795 131.295 20.965 ;
        RECT 131.125 15.355 131.295 15.525 ;
        RECT 131.125 9.915 131.295 10.085 ;
        RECT 131.585 58.875 131.755 59.045 ;
        RECT 131.585 53.435 131.755 53.605 ;
        RECT 131.585 47.995 131.755 48.165 ;
        RECT 131.585 42.555 131.755 42.725 ;
        RECT 131.585 37.115 131.755 37.285 ;
        RECT 131.585 31.675 131.755 31.845 ;
        RECT 131.585 26.235 131.755 26.405 ;
        RECT 131.585 20.795 131.755 20.965 ;
        RECT 131.585 15.355 131.755 15.525 ;
        RECT 131.585 9.915 131.755 10.085 ;
        RECT 132.045 58.875 132.215 59.045 ;
        RECT 132.045 53.435 132.215 53.605 ;
        RECT 132.045 47.995 132.215 48.165 ;
        RECT 132.045 42.555 132.215 42.725 ;
        RECT 132.045 37.115 132.215 37.285 ;
        RECT 132.045 31.675 132.215 31.845 ;
        RECT 132.045 26.235 132.215 26.405 ;
        RECT 132.045 20.795 132.215 20.965 ;
        RECT 132.045 15.355 132.215 15.525 ;
        RECT 132.045 9.915 132.215 10.085 ;
        RECT 132.505 58.875 132.675 59.045 ;
        RECT 132.505 53.435 132.675 53.605 ;
        RECT 132.505 47.995 132.675 48.165 ;
        RECT 132.505 42.555 132.675 42.725 ;
        RECT 132.505 37.115 132.675 37.285 ;
        RECT 132.505 31.675 132.675 31.845 ;
        RECT 132.505 26.235 132.675 26.405 ;
        RECT 132.505 20.795 132.675 20.965 ;
        RECT 132.505 15.355 132.675 15.525 ;
        RECT 132.505 9.915 132.675 10.085 ;
        RECT 132.965 58.875 133.135 59.045 ;
        RECT 132.965 53.435 133.135 53.605 ;
        RECT 132.965 47.995 133.135 48.165 ;
        RECT 132.965 42.555 133.135 42.725 ;
        RECT 132.965 37.115 133.135 37.285 ;
        RECT 132.965 31.675 133.135 31.845 ;
        RECT 132.965 26.235 133.135 26.405 ;
        RECT 132.965 20.795 133.135 20.965 ;
        RECT 132.965 15.355 133.135 15.525 ;
        RECT 132.965 9.915 133.135 10.085 ;
        RECT 133.425 58.875 133.595 59.045 ;
        RECT 133.425 53.435 133.595 53.605 ;
        RECT 133.425 47.995 133.595 48.165 ;
        RECT 133.425 42.555 133.595 42.725 ;
        RECT 133.425 37.115 133.595 37.285 ;
        RECT 133.425 31.675 133.595 31.845 ;
        RECT 133.425 26.235 133.595 26.405 ;
        RECT 133.425 20.795 133.595 20.965 ;
        RECT 133.425 15.355 133.595 15.525 ;
        RECT 133.425 9.915 133.595 10.085 ;
        RECT 133.885 58.875 134.055 59.045 ;
        RECT 133.885 53.435 134.055 53.605 ;
        RECT 133.885 47.995 134.055 48.165 ;
        RECT 133.885 42.555 134.055 42.725 ;
        RECT 133.885 37.115 134.055 37.285 ;
        RECT 133.885 31.675 134.055 31.845 ;
        RECT 133.885 26.235 134.055 26.405 ;
        RECT 133.885 20.795 134.055 20.965 ;
        RECT 133.885 15.355 134.055 15.525 ;
        RECT 133.885 9.915 134.055 10.085 ;
        RECT 134.345 58.875 134.515 59.045 ;
        RECT 134.345 53.435 134.515 53.605 ;
        RECT 134.345 47.995 134.515 48.165 ;
        RECT 134.345 42.555 134.515 42.725 ;
        RECT 134.345 37.115 134.515 37.285 ;
        RECT 134.345 31.675 134.515 31.845 ;
        RECT 134.345 26.235 134.515 26.405 ;
        RECT 134.345 20.795 134.515 20.965 ;
        RECT 134.345 15.355 134.515 15.525 ;
        RECT 134.345 9.915 134.515 10.085 ;
        RECT 134.805 58.875 134.975 59.045 ;
        RECT 134.805 53.435 134.975 53.605 ;
        RECT 134.805 47.995 134.975 48.165 ;
        RECT 134.805 42.555 134.975 42.725 ;
        RECT 134.805 37.115 134.975 37.285 ;
        RECT 134.805 31.675 134.975 31.845 ;
        RECT 134.805 26.235 134.975 26.405 ;
        RECT 134.805 20.795 134.975 20.965 ;
        RECT 134.805 15.355 134.975 15.525 ;
        RECT 134.805 9.915 134.975 10.085 ;
        RECT 135.265 58.875 135.435 59.045 ;
        RECT 135.265 53.435 135.435 53.605 ;
        RECT 135.265 47.995 135.435 48.165 ;
        RECT 135.265 42.555 135.435 42.725 ;
        RECT 135.265 37.115 135.435 37.285 ;
        RECT 135.265 31.675 135.435 31.845 ;
        RECT 135.265 26.235 135.435 26.405 ;
        RECT 135.265 20.795 135.435 20.965 ;
        RECT 135.265 15.355 135.435 15.525 ;
        RECT 135.265 9.915 135.435 10.085 ;
        RECT 135.725 58.875 135.895 59.045 ;
        RECT 135.725 53.435 135.895 53.605 ;
        RECT 135.725 47.995 135.895 48.165 ;
        RECT 135.725 42.555 135.895 42.725 ;
        RECT 135.725 37.115 135.895 37.285 ;
        RECT 135.725 31.675 135.895 31.845 ;
        RECT 135.725 26.235 135.895 26.405 ;
        RECT 135.725 20.795 135.895 20.965 ;
        RECT 135.725 15.355 135.895 15.525 ;
        RECT 135.725 9.915 135.895 10.085 ;
        RECT 136.185 58.875 136.355 59.045 ;
        RECT 136.185 53.435 136.355 53.605 ;
        RECT 136.185 47.995 136.355 48.165 ;
        RECT 136.185 42.555 136.355 42.725 ;
        RECT 136.185 37.115 136.355 37.285 ;
        RECT 136.185 31.675 136.355 31.845 ;
        RECT 136.185 26.235 136.355 26.405 ;
        RECT 136.185 20.795 136.355 20.965 ;
        RECT 136.185 15.355 136.355 15.525 ;
        RECT 136.185 9.915 136.355 10.085 ;
        RECT 136.645 58.875 136.815 59.045 ;
        RECT 136.645 53.435 136.815 53.605 ;
        RECT 136.645 47.995 136.815 48.165 ;
        RECT 136.645 42.555 136.815 42.725 ;
        RECT 136.645 37.115 136.815 37.285 ;
        RECT 136.645 31.675 136.815 31.845 ;
        RECT 136.645 26.235 136.815 26.405 ;
        RECT 136.645 20.795 136.815 20.965 ;
        RECT 136.645 15.355 136.815 15.525 ;
        RECT 136.645 9.915 136.815 10.085 ;
        RECT 137.105 58.875 137.275 59.045 ;
        RECT 137.105 53.435 137.275 53.605 ;
        RECT 137.105 47.995 137.275 48.165 ;
        RECT 137.105 42.555 137.275 42.725 ;
        RECT 137.105 37.115 137.275 37.285 ;
        RECT 137.105 31.675 137.275 31.845 ;
        RECT 137.105 26.235 137.275 26.405 ;
        RECT 137.105 20.795 137.275 20.965 ;
        RECT 137.105 15.355 137.275 15.525 ;
        RECT 137.105 9.915 137.275 10.085 ;
        RECT 137.565 58.875 137.735 59.045 ;
        RECT 137.565 53.435 137.735 53.605 ;
        RECT 137.565 47.995 137.735 48.165 ;
        RECT 137.565 42.555 137.735 42.725 ;
        RECT 137.565 37.115 137.735 37.285 ;
        RECT 137.565 31.675 137.735 31.845 ;
        RECT 137.565 26.235 137.735 26.405 ;
        RECT 137.565 20.795 137.735 20.965 ;
        RECT 137.565 15.355 137.735 15.525 ;
        RECT 137.565 9.915 137.735 10.085 ;
        RECT 138.025 58.875 138.195 59.045 ;
        RECT 138.025 53.435 138.195 53.605 ;
        RECT 138.025 47.995 138.195 48.165 ;
        RECT 138.025 42.555 138.195 42.725 ;
        RECT 138.025 37.115 138.195 37.285 ;
        RECT 138.025 31.675 138.195 31.845 ;
        RECT 138.025 26.235 138.195 26.405 ;
        RECT 138.025 20.795 138.195 20.965 ;
        RECT 138.025 15.355 138.195 15.525 ;
        RECT 138.025 9.915 138.195 10.085 ;
        RECT 138.485 58.875 138.655 59.045 ;
        RECT 138.485 53.435 138.655 53.605 ;
        RECT 138.485 47.995 138.655 48.165 ;
        RECT 138.485 42.555 138.655 42.725 ;
        RECT 138.485 37.115 138.655 37.285 ;
        RECT 138.485 31.675 138.655 31.845 ;
        RECT 138.485 26.235 138.655 26.405 ;
        RECT 138.485 20.795 138.655 20.965 ;
        RECT 138.485 15.355 138.655 15.525 ;
        RECT 138.485 9.915 138.655 10.085 ;
        RECT 138.945 58.875 139.115 59.045 ;
        RECT 138.945 53.435 139.115 53.605 ;
        RECT 138.945 47.995 139.115 48.165 ;
        RECT 138.945 42.555 139.115 42.725 ;
        RECT 138.945 37.115 139.115 37.285 ;
        RECT 138.945 31.675 139.115 31.845 ;
        RECT 138.945 26.235 139.115 26.405 ;
        RECT 138.945 20.795 139.115 20.965 ;
        RECT 138.945 15.355 139.115 15.525 ;
        RECT 138.945 9.915 139.115 10.085 ;
        RECT 139.405 58.875 139.575 59.045 ;
        RECT 139.405 53.435 139.575 53.605 ;
        RECT 139.405 47.995 139.575 48.165 ;
        RECT 139.405 42.555 139.575 42.725 ;
        RECT 139.405 37.115 139.575 37.285 ;
        RECT 139.405 31.675 139.575 31.845 ;
        RECT 139.405 26.235 139.575 26.405 ;
        RECT 139.405 20.795 139.575 20.965 ;
        RECT 139.405 15.355 139.575 15.525 ;
        RECT 139.405 9.915 139.575 10.085 ;
        RECT 139.865 58.875 140.035 59.045 ;
        RECT 139.865 53.435 140.035 53.605 ;
        RECT 139.865 47.995 140.035 48.165 ;
        RECT 139.865 42.555 140.035 42.725 ;
        RECT 139.865 37.115 140.035 37.285 ;
        RECT 139.865 31.675 140.035 31.845 ;
        RECT 139.865 26.235 140.035 26.405 ;
        RECT 139.865 20.795 140.035 20.965 ;
        RECT 139.865 15.355 140.035 15.525 ;
        RECT 139.865 9.915 140.035 10.085 ;
        RECT 140.325 58.875 140.495 59.045 ;
        RECT 140.325 53.435 140.495 53.605 ;
        RECT 140.325 47.995 140.495 48.165 ;
        RECT 140.325 42.555 140.495 42.725 ;
        RECT 140.325 37.115 140.495 37.285 ;
        RECT 140.325 31.675 140.495 31.845 ;
        RECT 140.325 26.235 140.495 26.405 ;
        RECT 140.325 20.795 140.495 20.965 ;
        RECT 140.325 15.355 140.495 15.525 ;
        RECT 140.325 9.915 140.495 10.085 ;
        RECT 140.785 58.875 140.955 59.045 ;
        RECT 140.785 53.435 140.955 53.605 ;
        RECT 140.785 47.995 140.955 48.165 ;
        RECT 140.785 42.555 140.955 42.725 ;
        RECT 140.785 37.115 140.955 37.285 ;
        RECT 140.785 31.675 140.955 31.845 ;
        RECT 140.785 26.235 140.955 26.405 ;
        RECT 140.785 20.795 140.955 20.965 ;
        RECT 140.785 15.355 140.955 15.525 ;
        RECT 140.785 9.915 140.955 10.085 ;
        RECT 141.245 58.875 141.415 59.045 ;
        RECT 141.245 53.435 141.415 53.605 ;
        RECT 141.245 47.995 141.415 48.165 ;
        RECT 141.245 42.555 141.415 42.725 ;
        RECT 141.245 37.115 141.415 37.285 ;
        RECT 141.245 31.675 141.415 31.845 ;
        RECT 141.245 26.235 141.415 26.405 ;
        RECT 141.245 20.795 141.415 20.965 ;
        RECT 141.245 15.355 141.415 15.525 ;
        RECT 141.245 9.915 141.415 10.085 ;
        RECT 141.705 58.875 141.875 59.045 ;
        RECT 141.705 53.435 141.875 53.605 ;
        RECT 141.705 47.995 141.875 48.165 ;
        RECT 141.705 42.555 141.875 42.725 ;
        RECT 141.705 37.115 141.875 37.285 ;
        RECT 141.705 31.675 141.875 31.845 ;
        RECT 141.705 26.235 141.875 26.405 ;
        RECT 141.705 20.795 141.875 20.965 ;
        RECT 141.705 15.355 141.875 15.525 ;
        RECT 141.705 9.915 141.875 10.085 ;
        RECT 142.165 58.875 142.335 59.045 ;
        RECT 142.165 53.435 142.335 53.605 ;
        RECT 142.165 47.995 142.335 48.165 ;
        RECT 142.165 42.555 142.335 42.725 ;
        RECT 142.165 37.115 142.335 37.285 ;
        RECT 142.165 31.675 142.335 31.845 ;
        RECT 142.165 26.235 142.335 26.405 ;
        RECT 142.165 20.795 142.335 20.965 ;
        RECT 142.165 15.355 142.335 15.525 ;
        RECT 142.165 9.915 142.335 10.085 ;
        RECT 142.625 58.875 142.795 59.045 ;
        RECT 142.625 53.435 142.795 53.605 ;
        RECT 142.625 47.995 142.795 48.165 ;
        RECT 142.625 42.555 142.795 42.725 ;
        RECT 142.625 37.115 142.795 37.285 ;
        RECT 142.625 31.675 142.795 31.845 ;
        RECT 142.625 26.235 142.795 26.405 ;
        RECT 142.625 20.795 142.795 20.965 ;
        RECT 142.625 15.355 142.795 15.525 ;
        RECT 142.625 9.915 142.795 10.085 ;
        RECT 143.085 58.875 143.255 59.045 ;
        RECT 143.085 53.435 143.255 53.605 ;
        RECT 143.085 47.995 143.255 48.165 ;
        RECT 143.085 42.555 143.255 42.725 ;
        RECT 143.085 37.115 143.255 37.285 ;
        RECT 143.085 31.675 143.255 31.845 ;
        RECT 143.085 26.235 143.255 26.405 ;
        RECT 143.085 20.795 143.255 20.965 ;
        RECT 143.085 15.355 143.255 15.525 ;
        RECT 143.085 9.915 143.255 10.085 ;
        RECT 143.545 58.875 143.715 59.045 ;
        RECT 143.545 53.435 143.715 53.605 ;
        RECT 143.545 47.995 143.715 48.165 ;
        RECT 143.545 42.555 143.715 42.725 ;
        RECT 143.545 37.115 143.715 37.285 ;
        RECT 143.545 31.675 143.715 31.845 ;
        RECT 143.545 26.235 143.715 26.405 ;
        RECT 143.545 20.795 143.715 20.965 ;
        RECT 143.545 15.355 143.715 15.525 ;
        RECT 143.545 9.915 143.715 10.085 ;
        RECT 144.005 58.875 144.175 59.045 ;
        RECT 144.005 53.435 144.175 53.605 ;
        RECT 144.005 47.995 144.175 48.165 ;
        RECT 144.005 42.555 144.175 42.725 ;
        RECT 144.005 37.115 144.175 37.285 ;
        RECT 144.005 31.675 144.175 31.845 ;
        RECT 144.005 26.235 144.175 26.405 ;
        RECT 144.005 20.795 144.175 20.965 ;
        RECT 144.005 15.355 144.175 15.525 ;
        RECT 144.005 9.915 144.175 10.085 ;
        RECT 144.465 58.875 144.635 59.045 ;
        RECT 144.465 53.435 144.635 53.605 ;
        RECT 144.465 47.995 144.635 48.165 ;
        RECT 144.465 42.555 144.635 42.725 ;
        RECT 144.465 37.115 144.635 37.285 ;
        RECT 144.465 31.675 144.635 31.845 ;
        RECT 144.465 26.235 144.635 26.405 ;
        RECT 144.465 20.795 144.635 20.965 ;
        RECT 144.465 15.355 144.635 15.525 ;
        RECT 144.465 9.915 144.635 10.085 ;
        RECT 144.925 58.875 145.095 59.045 ;
        RECT 144.925 53.435 145.095 53.605 ;
        RECT 144.925 47.995 145.095 48.165 ;
        RECT 144.925 42.555 145.095 42.725 ;
        RECT 144.925 37.115 145.095 37.285 ;
        RECT 144.925 31.675 145.095 31.845 ;
        RECT 144.925 26.235 145.095 26.405 ;
        RECT 144.925 20.795 145.095 20.965 ;
        RECT 144.925 15.355 145.095 15.525 ;
        RECT 144.925 9.915 145.095 10.085 ;
        RECT 145.385 58.875 145.555 59.045 ;
        RECT 145.385 53.435 145.555 53.605 ;
        RECT 145.385 47.995 145.555 48.165 ;
        RECT 145.385 42.555 145.555 42.725 ;
        RECT 145.385 37.115 145.555 37.285 ;
        RECT 145.385 31.675 145.555 31.845 ;
        RECT 145.385 26.235 145.555 26.405 ;
        RECT 145.385 20.795 145.555 20.965 ;
        RECT 145.385 15.355 145.555 15.525 ;
        RECT 145.385 9.915 145.555 10.085 ;
        RECT 145.845 58.875 146.015 59.045 ;
        RECT 145.845 53.435 146.015 53.605 ;
        RECT 145.845 47.995 146.015 48.165 ;
        RECT 145.845 42.555 146.015 42.725 ;
        RECT 145.845 37.115 146.015 37.285 ;
        RECT 145.845 31.675 146.015 31.845 ;
        RECT 145.845 26.235 146.015 26.405 ;
        RECT 145.845 20.795 146.015 20.965 ;
        RECT 145.845 15.355 146.015 15.525 ;
        RECT 145.845 9.915 146.015 10.085 ;
        RECT 146.305 58.875 146.475 59.045 ;
        RECT 146.305 53.435 146.475 53.605 ;
        RECT 146.305 47.995 146.475 48.165 ;
        RECT 146.305 42.555 146.475 42.725 ;
        RECT 146.305 37.115 146.475 37.285 ;
        RECT 146.305 31.675 146.475 31.845 ;
        RECT 146.305 26.235 146.475 26.405 ;
        RECT 146.305 20.795 146.475 20.965 ;
        RECT 146.305 15.355 146.475 15.525 ;
        RECT 146.305 9.915 146.475 10.085 ;
        RECT 146.765 58.875 146.935 59.045 ;
        RECT 146.765 53.435 146.935 53.605 ;
        RECT 146.765 47.995 146.935 48.165 ;
        RECT 146.765 42.555 146.935 42.725 ;
        RECT 146.765 37.115 146.935 37.285 ;
        RECT 146.765 31.675 146.935 31.845 ;
        RECT 146.765 26.235 146.935 26.405 ;
        RECT 146.765 20.795 146.935 20.965 ;
        RECT 146.765 15.355 146.935 15.525 ;
        RECT 146.765 9.915 146.935 10.085 ;
        RECT 147.225 58.875 147.395 59.045 ;
        RECT 147.225 53.435 147.395 53.605 ;
        RECT 147.225 47.995 147.395 48.165 ;
        RECT 147.225 42.555 147.395 42.725 ;
        RECT 147.225 37.115 147.395 37.285 ;
        RECT 147.225 31.675 147.395 31.845 ;
        RECT 147.225 26.235 147.395 26.405 ;
        RECT 147.225 20.795 147.395 20.965 ;
        RECT 147.225 15.355 147.395 15.525 ;
        RECT 147.225 9.915 147.395 10.085 ;
        RECT 147.685 58.875 147.855 59.045 ;
        RECT 147.685 53.435 147.855 53.605 ;
        RECT 147.685 47.995 147.855 48.165 ;
        RECT 147.685 42.555 147.855 42.725 ;
        RECT 147.685 37.115 147.855 37.285 ;
        RECT 147.685 31.675 147.855 31.845 ;
        RECT 147.685 26.235 147.855 26.405 ;
        RECT 147.685 20.795 147.855 20.965 ;
        RECT 147.685 15.355 147.855 15.525 ;
        RECT 147.685 9.915 147.855 10.085 ;
        RECT 56.145 58.875 56.315 59.045 ;
        RECT 56.145 53.435 56.315 53.605 ;
        RECT 56.145 47.995 56.315 48.165 ;
        RECT 56.145 42.555 56.315 42.725 ;
        RECT 56.145 37.115 56.315 37.285 ;
        RECT 56.145 31.675 56.315 31.845 ;
        RECT 56.145 26.235 56.315 26.405 ;
        RECT 56.145 20.795 56.315 20.965 ;
        RECT 56.145 15.355 56.315 15.525 ;
        RECT 56.145 9.915 56.315 10.085 ;
        RECT 56.605 58.875 56.775 59.045 ;
        RECT 56.605 53.435 56.775 53.605 ;
        RECT 56.605 47.995 56.775 48.165 ;
        RECT 56.605 42.555 56.775 42.725 ;
        RECT 56.605 37.115 56.775 37.285 ;
        RECT 56.605 31.675 56.775 31.845 ;
        RECT 56.605 26.235 56.775 26.405 ;
        RECT 56.605 20.795 56.775 20.965 ;
        RECT 56.605 15.355 56.775 15.525 ;
        RECT 56.605 9.915 56.775 10.085 ;
        RECT 57.065 58.875 57.235 59.045 ;
        RECT 57.065 53.435 57.235 53.605 ;
        RECT 57.065 47.995 57.235 48.165 ;
        RECT 57.065 42.555 57.235 42.725 ;
        RECT 57.065 37.115 57.235 37.285 ;
        RECT 57.065 31.675 57.235 31.845 ;
        RECT 57.065 26.235 57.235 26.405 ;
        RECT 57.065 20.795 57.235 20.965 ;
        RECT 57.065 15.355 57.235 15.525 ;
        RECT 57.065 9.915 57.235 10.085 ;
        RECT 57.525 58.875 57.695 59.045 ;
        RECT 57.525 53.435 57.695 53.605 ;
        RECT 57.525 47.995 57.695 48.165 ;
        RECT 57.525 42.555 57.695 42.725 ;
        RECT 57.525 37.115 57.695 37.285 ;
        RECT 57.525 31.675 57.695 31.845 ;
        RECT 57.525 26.235 57.695 26.405 ;
        RECT 57.525 20.795 57.695 20.965 ;
        RECT 57.525 15.355 57.695 15.525 ;
        RECT 57.525 9.915 57.695 10.085 ;
        RECT 57.985 58.875 58.155 59.045 ;
        RECT 57.985 53.435 58.155 53.605 ;
        RECT 57.985 47.995 58.155 48.165 ;
        RECT 57.985 42.555 58.155 42.725 ;
        RECT 57.985 37.115 58.155 37.285 ;
        RECT 57.985 31.675 58.155 31.845 ;
        RECT 57.985 26.235 58.155 26.405 ;
        RECT 57.985 20.795 58.155 20.965 ;
        RECT 57.985 15.355 58.155 15.525 ;
        RECT 57.985 9.915 58.155 10.085 ;
        RECT 58.445 58.875 58.615 59.045 ;
        RECT 58.445 53.435 58.615 53.605 ;
        RECT 58.445 47.995 58.615 48.165 ;
        RECT 58.445 42.555 58.615 42.725 ;
        RECT 58.445 37.115 58.615 37.285 ;
        RECT 58.445 31.675 58.615 31.845 ;
        RECT 58.445 26.235 58.615 26.405 ;
        RECT 58.445 20.795 58.615 20.965 ;
        RECT 58.445 15.355 58.615 15.525 ;
        RECT 58.445 9.915 58.615 10.085 ;
        RECT 58.905 58.875 59.075 59.045 ;
        RECT 58.905 53.435 59.075 53.605 ;
        RECT 58.905 47.995 59.075 48.165 ;
        RECT 58.905 42.555 59.075 42.725 ;
        RECT 58.905 37.115 59.075 37.285 ;
        RECT 58.905 31.675 59.075 31.845 ;
        RECT 58.905 26.235 59.075 26.405 ;
        RECT 58.905 20.795 59.075 20.965 ;
        RECT 58.905 15.355 59.075 15.525 ;
        RECT 58.905 9.915 59.075 10.085 ;
        RECT 59.365 58.875 59.535 59.045 ;
        RECT 59.365 53.435 59.535 53.605 ;
        RECT 59.365 47.995 59.535 48.165 ;
        RECT 59.365 42.555 59.535 42.725 ;
        RECT 59.365 37.115 59.535 37.285 ;
        RECT 59.365 31.675 59.535 31.845 ;
        RECT 59.365 26.235 59.535 26.405 ;
        RECT 59.365 20.795 59.535 20.965 ;
        RECT 59.365 15.355 59.535 15.525 ;
        RECT 59.365 9.915 59.535 10.085 ;
        RECT 59.825 58.875 59.995 59.045 ;
        RECT 59.825 53.435 59.995 53.605 ;
        RECT 59.825 47.995 59.995 48.165 ;
        RECT 59.825 42.555 59.995 42.725 ;
        RECT 59.825 37.115 59.995 37.285 ;
        RECT 59.825 31.675 59.995 31.845 ;
        RECT 59.825 26.235 59.995 26.405 ;
        RECT 59.825 20.795 59.995 20.965 ;
        RECT 59.825 15.355 59.995 15.525 ;
        RECT 59.825 9.915 59.995 10.085 ;
        RECT 60.285 58.875 60.455 59.045 ;
        RECT 60.285 53.435 60.455 53.605 ;
        RECT 60.285 47.995 60.455 48.165 ;
        RECT 60.285 42.555 60.455 42.725 ;
        RECT 60.285 37.115 60.455 37.285 ;
        RECT 60.285 31.675 60.455 31.845 ;
        RECT 60.285 26.235 60.455 26.405 ;
        RECT 60.285 20.795 60.455 20.965 ;
        RECT 60.285 15.355 60.455 15.525 ;
        RECT 60.285 9.915 60.455 10.085 ;
        RECT 60.745 58.875 60.915 59.045 ;
        RECT 60.745 53.435 60.915 53.605 ;
        RECT 60.745 47.995 60.915 48.165 ;
        RECT 60.745 42.555 60.915 42.725 ;
        RECT 60.745 37.115 60.915 37.285 ;
        RECT 60.745 31.675 60.915 31.845 ;
        RECT 60.745 26.235 60.915 26.405 ;
        RECT 60.745 20.795 60.915 20.965 ;
        RECT 60.745 15.355 60.915 15.525 ;
        RECT 60.745 9.915 60.915 10.085 ;
        RECT 61.205 58.875 61.375 59.045 ;
        RECT 61.205 53.435 61.375 53.605 ;
        RECT 61.205 47.995 61.375 48.165 ;
        RECT 61.205 42.555 61.375 42.725 ;
        RECT 61.205 37.115 61.375 37.285 ;
        RECT 61.205 31.675 61.375 31.845 ;
        RECT 61.205 26.235 61.375 26.405 ;
        RECT 61.205 20.795 61.375 20.965 ;
        RECT 61.205 15.355 61.375 15.525 ;
        RECT 61.205 9.915 61.375 10.085 ;
        RECT 61.665 58.875 61.835 59.045 ;
        RECT 61.665 53.435 61.835 53.605 ;
        RECT 61.665 47.995 61.835 48.165 ;
        RECT 61.665 42.555 61.835 42.725 ;
        RECT 61.665 37.115 61.835 37.285 ;
        RECT 61.665 31.675 61.835 31.845 ;
        RECT 61.665 26.235 61.835 26.405 ;
        RECT 61.665 20.795 61.835 20.965 ;
        RECT 61.665 15.355 61.835 15.525 ;
        RECT 61.665 9.915 61.835 10.085 ;
        RECT 62.125 58.875 62.295 59.045 ;
        RECT 62.125 53.435 62.295 53.605 ;
        RECT 62.125 47.995 62.295 48.165 ;
        RECT 62.125 42.555 62.295 42.725 ;
        RECT 62.125 37.115 62.295 37.285 ;
        RECT 62.125 31.675 62.295 31.845 ;
        RECT 62.125 26.235 62.295 26.405 ;
        RECT 62.125 20.795 62.295 20.965 ;
        RECT 62.125 15.355 62.295 15.525 ;
        RECT 62.125 9.915 62.295 10.085 ;
        RECT 62.585 58.875 62.755 59.045 ;
        RECT 62.585 53.435 62.755 53.605 ;
        RECT 62.585 47.995 62.755 48.165 ;
        RECT 62.585 42.555 62.755 42.725 ;
        RECT 62.585 37.115 62.755 37.285 ;
        RECT 62.585 31.675 62.755 31.845 ;
        RECT 62.585 26.235 62.755 26.405 ;
        RECT 62.585 20.795 62.755 20.965 ;
        RECT 62.585 15.355 62.755 15.525 ;
        RECT 62.585 9.915 62.755 10.085 ;
        RECT 63.045 58.875 63.215 59.045 ;
        RECT 63.045 53.435 63.215 53.605 ;
        RECT 63.045 47.995 63.215 48.165 ;
        RECT 63.045 42.555 63.215 42.725 ;
        RECT 63.045 37.115 63.215 37.285 ;
        RECT 63.045 31.675 63.215 31.845 ;
        RECT 63.045 26.235 63.215 26.405 ;
        RECT 63.045 20.795 63.215 20.965 ;
        RECT 63.045 15.355 63.215 15.525 ;
        RECT 63.045 9.915 63.215 10.085 ;
        RECT 63.505 58.875 63.675 59.045 ;
        RECT 63.505 53.435 63.675 53.605 ;
        RECT 63.505 47.995 63.675 48.165 ;
        RECT 63.505 42.555 63.675 42.725 ;
        RECT 63.505 37.115 63.675 37.285 ;
        RECT 63.505 31.675 63.675 31.845 ;
        RECT 63.505 26.235 63.675 26.405 ;
        RECT 63.505 20.795 63.675 20.965 ;
        RECT 63.505 15.355 63.675 15.525 ;
        RECT 63.505 9.915 63.675 10.085 ;
        RECT 63.965 58.875 64.135 59.045 ;
        RECT 63.965 53.435 64.135 53.605 ;
        RECT 63.965 47.995 64.135 48.165 ;
        RECT 63.965 42.555 64.135 42.725 ;
        RECT 63.965 37.115 64.135 37.285 ;
        RECT 63.965 31.675 64.135 31.845 ;
        RECT 63.965 26.235 64.135 26.405 ;
        RECT 63.965 20.795 64.135 20.965 ;
        RECT 63.965 15.355 64.135 15.525 ;
        RECT 63.965 9.915 64.135 10.085 ;
        RECT 64.425 58.875 64.595 59.045 ;
        RECT 64.425 53.435 64.595 53.605 ;
        RECT 64.425 47.995 64.595 48.165 ;
        RECT 64.425 42.555 64.595 42.725 ;
        RECT 64.425 37.115 64.595 37.285 ;
        RECT 64.425 31.675 64.595 31.845 ;
        RECT 64.425 26.235 64.595 26.405 ;
        RECT 64.425 20.795 64.595 20.965 ;
        RECT 64.425 15.355 64.595 15.525 ;
        RECT 64.425 9.915 64.595 10.085 ;
        RECT 64.885 58.875 65.055 59.045 ;
        RECT 64.885 53.435 65.055 53.605 ;
        RECT 64.885 47.995 65.055 48.165 ;
        RECT 64.885 42.555 65.055 42.725 ;
        RECT 64.885 37.115 65.055 37.285 ;
        RECT 64.885 31.675 65.055 31.845 ;
        RECT 64.885 26.235 65.055 26.405 ;
        RECT 64.885 20.795 65.055 20.965 ;
        RECT 64.885 15.355 65.055 15.525 ;
        RECT 64.885 9.915 65.055 10.085 ;
        RECT 65.345 58.875 65.515 59.045 ;
        RECT 65.345 53.435 65.515 53.605 ;
        RECT 65.345 47.995 65.515 48.165 ;
        RECT 65.345 42.555 65.515 42.725 ;
        RECT 65.345 37.115 65.515 37.285 ;
        RECT 65.345 31.675 65.515 31.845 ;
        RECT 65.345 26.235 65.515 26.405 ;
        RECT 65.345 20.795 65.515 20.965 ;
        RECT 65.345 15.355 65.515 15.525 ;
        RECT 65.345 9.915 65.515 10.085 ;
        RECT 65.805 58.875 65.975 59.045 ;
        RECT 65.805 53.435 65.975 53.605 ;
        RECT 65.805 47.995 65.975 48.165 ;
        RECT 65.805 42.555 65.975 42.725 ;
        RECT 65.805 37.115 65.975 37.285 ;
        RECT 65.805 31.675 65.975 31.845 ;
        RECT 65.805 26.235 65.975 26.405 ;
        RECT 65.805 20.795 65.975 20.965 ;
        RECT 65.805 15.355 65.975 15.525 ;
        RECT 65.805 9.915 65.975 10.085 ;
        RECT 66.265 58.875 66.435 59.045 ;
        RECT 66.265 53.435 66.435 53.605 ;
        RECT 66.265 47.995 66.435 48.165 ;
        RECT 66.265 42.555 66.435 42.725 ;
        RECT 66.265 37.115 66.435 37.285 ;
        RECT 66.265 31.675 66.435 31.845 ;
        RECT 66.265 26.235 66.435 26.405 ;
        RECT 66.265 20.795 66.435 20.965 ;
        RECT 66.265 15.355 66.435 15.525 ;
        RECT 66.265 9.915 66.435 10.085 ;
        RECT 66.725 58.875 66.895 59.045 ;
        RECT 66.725 53.435 66.895 53.605 ;
        RECT 66.725 47.995 66.895 48.165 ;
        RECT 66.725 42.555 66.895 42.725 ;
        RECT 66.725 37.115 66.895 37.285 ;
        RECT 66.725 31.675 66.895 31.845 ;
        RECT 66.725 26.235 66.895 26.405 ;
        RECT 66.725 20.795 66.895 20.965 ;
        RECT 66.725 15.355 66.895 15.525 ;
        RECT 66.725 9.915 66.895 10.085 ;
        RECT 67.185 58.875 67.355 59.045 ;
        RECT 67.185 53.435 67.355 53.605 ;
        RECT 67.185 47.995 67.355 48.165 ;
        RECT 67.185 42.555 67.355 42.725 ;
        RECT 67.185 37.115 67.355 37.285 ;
        RECT 67.185 31.675 67.355 31.845 ;
        RECT 67.185 26.235 67.355 26.405 ;
        RECT 67.185 20.795 67.355 20.965 ;
        RECT 67.185 15.355 67.355 15.525 ;
        RECT 67.185 9.915 67.355 10.085 ;
        RECT 67.645 58.875 67.815 59.045 ;
        RECT 67.645 53.435 67.815 53.605 ;
        RECT 67.645 47.995 67.815 48.165 ;
        RECT 67.645 42.555 67.815 42.725 ;
        RECT 67.645 37.115 67.815 37.285 ;
        RECT 67.645 31.675 67.815 31.845 ;
        RECT 67.645 26.235 67.815 26.405 ;
        RECT 67.645 20.795 67.815 20.965 ;
        RECT 67.645 15.355 67.815 15.525 ;
        RECT 67.645 9.915 67.815 10.085 ;
        RECT 68.105 58.875 68.275 59.045 ;
        RECT 68.105 53.435 68.275 53.605 ;
        RECT 68.105 47.995 68.275 48.165 ;
        RECT 68.105 42.555 68.275 42.725 ;
        RECT 68.105 37.115 68.275 37.285 ;
        RECT 68.105 31.675 68.275 31.845 ;
        RECT 68.105 26.235 68.275 26.405 ;
        RECT 68.105 20.795 68.275 20.965 ;
        RECT 68.105 15.355 68.275 15.525 ;
        RECT 68.105 9.915 68.275 10.085 ;
        RECT 68.565 58.875 68.735 59.045 ;
        RECT 68.565 53.435 68.735 53.605 ;
        RECT 68.565 47.995 68.735 48.165 ;
        RECT 68.565 42.555 68.735 42.725 ;
        RECT 68.565 37.115 68.735 37.285 ;
        RECT 68.565 31.675 68.735 31.845 ;
        RECT 68.565 26.235 68.735 26.405 ;
        RECT 68.565 20.795 68.735 20.965 ;
        RECT 68.565 15.355 68.735 15.525 ;
        RECT 68.565 9.915 68.735 10.085 ;
        RECT 69.025 58.875 69.195 59.045 ;
        RECT 69.025 53.435 69.195 53.605 ;
        RECT 69.025 47.995 69.195 48.165 ;
        RECT 69.025 42.555 69.195 42.725 ;
        RECT 69.025 37.115 69.195 37.285 ;
        RECT 69.025 31.675 69.195 31.845 ;
        RECT 69.025 26.235 69.195 26.405 ;
        RECT 69.025 20.795 69.195 20.965 ;
        RECT 69.025 15.355 69.195 15.525 ;
        RECT 69.025 9.915 69.195 10.085 ;
        RECT 69.485 58.875 69.655 59.045 ;
        RECT 69.485 53.435 69.655 53.605 ;
        RECT 69.485 47.995 69.655 48.165 ;
        RECT 69.485 42.555 69.655 42.725 ;
        RECT 69.485 37.115 69.655 37.285 ;
        RECT 69.485 31.675 69.655 31.845 ;
        RECT 69.485 26.235 69.655 26.405 ;
        RECT 69.485 20.795 69.655 20.965 ;
        RECT 69.485 15.355 69.655 15.525 ;
        RECT 69.485 9.915 69.655 10.085 ;
        RECT 69.945 58.875 70.115 59.045 ;
        RECT 69.945 53.435 70.115 53.605 ;
        RECT 69.945 47.995 70.115 48.165 ;
        RECT 69.945 42.555 70.115 42.725 ;
        RECT 69.945 37.115 70.115 37.285 ;
        RECT 69.945 31.675 70.115 31.845 ;
        RECT 69.945 26.235 70.115 26.405 ;
        RECT 69.945 20.795 70.115 20.965 ;
        RECT 69.945 15.355 70.115 15.525 ;
        RECT 69.945 9.915 70.115 10.085 ;
        RECT 70.405 58.875 70.575 59.045 ;
        RECT 70.405 53.435 70.575 53.605 ;
        RECT 70.405 47.995 70.575 48.165 ;
        RECT 70.405 42.555 70.575 42.725 ;
        RECT 70.405 37.115 70.575 37.285 ;
        RECT 70.405 31.675 70.575 31.845 ;
        RECT 70.405 26.235 70.575 26.405 ;
        RECT 70.405 20.795 70.575 20.965 ;
        RECT 70.405 15.355 70.575 15.525 ;
        RECT 70.405 9.915 70.575 10.085 ;
        RECT 70.865 58.875 71.035 59.045 ;
        RECT 70.865 53.435 71.035 53.605 ;
        RECT 70.865 47.995 71.035 48.165 ;
        RECT 70.865 42.555 71.035 42.725 ;
        RECT 70.865 37.115 71.035 37.285 ;
        RECT 70.865 31.675 71.035 31.845 ;
        RECT 70.865 26.235 71.035 26.405 ;
        RECT 70.865 20.795 71.035 20.965 ;
        RECT 70.865 15.355 71.035 15.525 ;
        RECT 70.865 9.915 71.035 10.085 ;
        RECT 71.325 58.875 71.495 59.045 ;
        RECT 71.325 53.435 71.495 53.605 ;
        RECT 71.325 47.995 71.495 48.165 ;
        RECT 71.325 42.555 71.495 42.725 ;
        RECT 71.325 37.115 71.495 37.285 ;
        RECT 71.325 31.675 71.495 31.845 ;
        RECT 71.325 26.235 71.495 26.405 ;
        RECT 71.325 20.795 71.495 20.965 ;
        RECT 71.325 15.355 71.495 15.525 ;
        RECT 71.325 9.915 71.495 10.085 ;
        RECT 71.785 58.875 71.955 59.045 ;
        RECT 71.785 53.435 71.955 53.605 ;
        RECT 71.785 47.995 71.955 48.165 ;
        RECT 71.785 42.555 71.955 42.725 ;
        RECT 71.785 37.115 71.955 37.285 ;
        RECT 71.785 31.675 71.955 31.845 ;
        RECT 71.785 26.235 71.955 26.405 ;
        RECT 71.785 20.795 71.955 20.965 ;
        RECT 71.785 15.355 71.955 15.525 ;
        RECT 71.785 9.915 71.955 10.085 ;
        RECT 72.245 58.875 72.415 59.045 ;
        RECT 72.245 53.435 72.415 53.605 ;
        RECT 72.245 47.995 72.415 48.165 ;
        RECT 72.245 42.555 72.415 42.725 ;
        RECT 72.245 37.115 72.415 37.285 ;
        RECT 72.245 31.675 72.415 31.845 ;
        RECT 72.245 26.235 72.415 26.405 ;
        RECT 72.245 20.795 72.415 20.965 ;
        RECT 72.245 15.355 72.415 15.525 ;
        RECT 72.245 9.915 72.415 10.085 ;
        RECT 72.705 58.875 72.875 59.045 ;
        RECT 72.705 53.435 72.875 53.605 ;
        RECT 72.705 47.995 72.875 48.165 ;
        RECT 72.705 42.555 72.875 42.725 ;
        RECT 72.705 37.115 72.875 37.285 ;
        RECT 72.705 31.675 72.875 31.845 ;
        RECT 72.705 26.235 72.875 26.405 ;
        RECT 72.705 20.795 72.875 20.965 ;
        RECT 72.705 15.355 72.875 15.525 ;
        RECT 72.705 9.915 72.875 10.085 ;
        RECT 73.165 58.875 73.335 59.045 ;
        RECT 73.165 53.435 73.335 53.605 ;
        RECT 73.165 47.995 73.335 48.165 ;
        RECT 73.165 42.555 73.335 42.725 ;
        RECT 73.165 37.115 73.335 37.285 ;
        RECT 73.165 31.675 73.335 31.845 ;
        RECT 73.165 26.235 73.335 26.405 ;
        RECT 73.165 20.795 73.335 20.965 ;
        RECT 73.165 15.355 73.335 15.525 ;
        RECT 73.165 9.915 73.335 10.085 ;
        RECT 73.625 58.875 73.795 59.045 ;
        RECT 73.625 53.435 73.795 53.605 ;
        RECT 73.625 47.995 73.795 48.165 ;
        RECT 73.625 42.555 73.795 42.725 ;
        RECT 73.625 37.115 73.795 37.285 ;
        RECT 73.625 31.675 73.795 31.845 ;
        RECT 73.625 26.235 73.795 26.405 ;
        RECT 73.625 20.795 73.795 20.965 ;
        RECT 73.625 15.355 73.795 15.525 ;
        RECT 73.625 9.915 73.795 10.085 ;
        RECT 74.085 58.875 74.255 59.045 ;
        RECT 74.085 53.435 74.255 53.605 ;
        RECT 74.085 47.995 74.255 48.165 ;
        RECT 74.085 42.555 74.255 42.725 ;
        RECT 74.085 37.115 74.255 37.285 ;
        RECT 74.085 31.675 74.255 31.845 ;
        RECT 74.085 26.235 74.255 26.405 ;
        RECT 74.085 20.795 74.255 20.965 ;
        RECT 74.085 15.355 74.255 15.525 ;
        RECT 74.085 9.915 74.255 10.085 ;
        RECT 74.545 58.875 74.715 59.045 ;
        RECT 74.545 53.435 74.715 53.605 ;
        RECT 74.545 47.995 74.715 48.165 ;
        RECT 74.545 42.555 74.715 42.725 ;
        RECT 74.545 37.115 74.715 37.285 ;
        RECT 74.545 31.675 74.715 31.845 ;
        RECT 74.545 26.235 74.715 26.405 ;
        RECT 74.545 20.795 74.715 20.965 ;
        RECT 74.545 15.355 74.715 15.525 ;
        RECT 74.545 9.915 74.715 10.085 ;
        RECT 75.005 58.875 75.175 59.045 ;
        RECT 75.005 53.435 75.175 53.605 ;
        RECT 75.005 47.995 75.175 48.165 ;
        RECT 75.005 42.555 75.175 42.725 ;
        RECT 75.005 37.115 75.175 37.285 ;
        RECT 75.005 31.675 75.175 31.845 ;
        RECT 75.005 26.235 75.175 26.405 ;
        RECT 75.005 20.795 75.175 20.965 ;
        RECT 75.005 15.355 75.175 15.525 ;
        RECT 75.005 9.915 75.175 10.085 ;
        RECT 75.465 58.875 75.635 59.045 ;
        RECT 75.465 53.435 75.635 53.605 ;
        RECT 75.465 47.995 75.635 48.165 ;
        RECT 75.465 42.555 75.635 42.725 ;
        RECT 75.465 37.115 75.635 37.285 ;
        RECT 75.465 31.675 75.635 31.845 ;
        RECT 75.465 26.235 75.635 26.405 ;
        RECT 75.465 20.795 75.635 20.965 ;
        RECT 75.465 15.355 75.635 15.525 ;
        RECT 75.465 9.915 75.635 10.085 ;
        RECT 75.925 58.875 76.095 59.045 ;
        RECT 75.925 53.435 76.095 53.605 ;
        RECT 75.925 47.995 76.095 48.165 ;
        RECT 75.925 42.555 76.095 42.725 ;
        RECT 75.925 37.115 76.095 37.285 ;
        RECT 75.925 31.675 76.095 31.845 ;
        RECT 75.925 26.235 76.095 26.405 ;
        RECT 75.925 20.795 76.095 20.965 ;
        RECT 75.925 15.355 76.095 15.525 ;
        RECT 75.925 9.915 76.095 10.085 ;
        RECT 76.385 58.875 76.555 59.045 ;
        RECT 76.385 53.435 76.555 53.605 ;
        RECT 76.385 47.995 76.555 48.165 ;
        RECT 76.385 42.555 76.555 42.725 ;
        RECT 76.385 37.115 76.555 37.285 ;
        RECT 76.385 31.675 76.555 31.845 ;
        RECT 76.385 26.235 76.555 26.405 ;
        RECT 76.385 20.795 76.555 20.965 ;
        RECT 76.385 15.355 76.555 15.525 ;
        RECT 76.385 9.915 76.555 10.085 ;
        RECT 76.845 58.875 77.015 59.045 ;
        RECT 76.845 53.435 77.015 53.605 ;
        RECT 76.845 47.995 77.015 48.165 ;
        RECT 76.845 42.555 77.015 42.725 ;
        RECT 76.845 37.115 77.015 37.285 ;
        RECT 76.845 31.675 77.015 31.845 ;
        RECT 76.845 26.235 77.015 26.405 ;
        RECT 76.845 20.795 77.015 20.965 ;
        RECT 76.845 15.355 77.015 15.525 ;
        RECT 76.845 9.915 77.015 10.085 ;
        RECT 77.305 58.875 77.475 59.045 ;
        RECT 77.305 53.435 77.475 53.605 ;
        RECT 77.305 47.995 77.475 48.165 ;
        RECT 77.305 42.555 77.475 42.725 ;
        RECT 77.305 37.115 77.475 37.285 ;
        RECT 77.305 31.675 77.475 31.845 ;
        RECT 77.305 26.235 77.475 26.405 ;
        RECT 77.305 20.795 77.475 20.965 ;
        RECT 77.305 15.355 77.475 15.525 ;
        RECT 77.305 9.915 77.475 10.085 ;
        RECT 77.765 58.875 77.935 59.045 ;
        RECT 77.765 53.435 77.935 53.605 ;
        RECT 77.765 47.995 77.935 48.165 ;
        RECT 77.765 42.555 77.935 42.725 ;
        RECT 77.765 37.115 77.935 37.285 ;
        RECT 77.765 31.675 77.935 31.845 ;
        RECT 77.765 26.235 77.935 26.405 ;
        RECT 77.765 20.795 77.935 20.965 ;
        RECT 77.765 15.355 77.935 15.525 ;
        RECT 77.765 9.915 77.935 10.085 ;
        RECT 78.225 58.875 78.395 59.045 ;
        RECT 78.225 53.435 78.395 53.605 ;
        RECT 78.225 47.995 78.395 48.165 ;
        RECT 78.225 42.555 78.395 42.725 ;
        RECT 78.225 37.115 78.395 37.285 ;
        RECT 78.225 31.675 78.395 31.845 ;
        RECT 78.225 26.235 78.395 26.405 ;
        RECT 78.225 20.795 78.395 20.965 ;
        RECT 78.225 15.355 78.395 15.525 ;
        RECT 78.225 9.915 78.395 10.085 ;
        RECT 78.685 58.875 78.855 59.045 ;
        RECT 78.685 53.435 78.855 53.605 ;
        RECT 78.685 47.995 78.855 48.165 ;
        RECT 78.685 42.555 78.855 42.725 ;
        RECT 78.685 37.115 78.855 37.285 ;
        RECT 78.685 31.675 78.855 31.845 ;
        RECT 78.685 26.235 78.855 26.405 ;
        RECT 78.685 20.795 78.855 20.965 ;
        RECT 78.685 15.355 78.855 15.525 ;
        RECT 78.685 9.915 78.855 10.085 ;
        RECT 79.145 58.875 79.315 59.045 ;
        RECT 79.145 53.435 79.315 53.605 ;
        RECT 79.145 47.995 79.315 48.165 ;
        RECT 79.145 42.555 79.315 42.725 ;
        RECT 79.145 37.115 79.315 37.285 ;
        RECT 79.145 31.675 79.315 31.845 ;
        RECT 79.145 26.235 79.315 26.405 ;
        RECT 79.145 20.795 79.315 20.965 ;
        RECT 79.145 15.355 79.315 15.525 ;
        RECT 79.145 9.915 79.315 10.085 ;
        RECT 79.605 58.875 79.775 59.045 ;
        RECT 79.605 53.435 79.775 53.605 ;
        RECT 79.605 47.995 79.775 48.165 ;
        RECT 79.605 42.555 79.775 42.725 ;
        RECT 79.605 37.115 79.775 37.285 ;
        RECT 79.605 31.675 79.775 31.845 ;
        RECT 79.605 26.235 79.775 26.405 ;
        RECT 79.605 20.795 79.775 20.965 ;
        RECT 79.605 15.355 79.775 15.525 ;
        RECT 79.605 9.915 79.775 10.085 ;
        RECT 80.065 58.875 80.235 59.045 ;
        RECT 80.065 53.435 80.235 53.605 ;
        RECT 80.065 47.995 80.235 48.165 ;
        RECT 80.065 42.555 80.235 42.725 ;
        RECT 80.065 37.115 80.235 37.285 ;
        RECT 80.065 31.675 80.235 31.845 ;
        RECT 80.065 26.235 80.235 26.405 ;
        RECT 80.065 20.795 80.235 20.965 ;
        RECT 80.065 15.355 80.235 15.525 ;
        RECT 80.065 9.915 80.235 10.085 ;
        RECT 80.525 58.875 80.695 59.045 ;
        RECT 80.525 53.435 80.695 53.605 ;
        RECT 80.525 47.995 80.695 48.165 ;
        RECT 80.525 42.555 80.695 42.725 ;
        RECT 80.525 37.115 80.695 37.285 ;
        RECT 80.525 31.675 80.695 31.845 ;
        RECT 80.525 26.235 80.695 26.405 ;
        RECT 80.525 20.795 80.695 20.965 ;
        RECT 80.525 15.355 80.695 15.525 ;
        RECT 80.525 9.915 80.695 10.085 ;
        RECT 80.985 58.875 81.155 59.045 ;
        RECT 80.985 53.435 81.155 53.605 ;
        RECT 80.985 47.995 81.155 48.165 ;
        RECT 80.985 42.555 81.155 42.725 ;
        RECT 80.985 37.115 81.155 37.285 ;
        RECT 80.985 31.675 81.155 31.845 ;
        RECT 80.985 26.235 81.155 26.405 ;
        RECT 80.985 20.795 81.155 20.965 ;
        RECT 80.985 15.355 81.155 15.525 ;
        RECT 80.985 9.915 81.155 10.085 ;
        RECT 81.445 58.875 81.615 59.045 ;
        RECT 81.445 53.435 81.615 53.605 ;
        RECT 81.445 47.995 81.615 48.165 ;
        RECT 81.445 42.555 81.615 42.725 ;
        RECT 81.445 37.115 81.615 37.285 ;
        RECT 81.445 31.675 81.615 31.845 ;
        RECT 81.445 26.235 81.615 26.405 ;
        RECT 81.445 20.795 81.615 20.965 ;
        RECT 81.445 15.355 81.615 15.525 ;
        RECT 81.445 9.915 81.615 10.085 ;
        RECT 81.905 58.875 82.075 59.045 ;
        RECT 81.905 53.435 82.075 53.605 ;
        RECT 81.905 47.995 82.075 48.165 ;
        RECT 81.905 42.555 82.075 42.725 ;
        RECT 81.905 37.115 82.075 37.285 ;
        RECT 81.905 31.675 82.075 31.845 ;
        RECT 81.905 26.235 82.075 26.405 ;
        RECT 81.905 20.795 82.075 20.965 ;
        RECT 81.905 15.355 82.075 15.525 ;
        RECT 81.905 9.915 82.075 10.085 ;
        RECT 82.365 58.875 82.535 59.045 ;
        RECT 82.365 53.435 82.535 53.605 ;
        RECT 82.365 47.995 82.535 48.165 ;
        RECT 82.365 42.555 82.535 42.725 ;
        RECT 82.365 37.115 82.535 37.285 ;
        RECT 82.365 31.675 82.535 31.845 ;
        RECT 82.365 26.235 82.535 26.405 ;
        RECT 82.365 20.795 82.535 20.965 ;
        RECT 82.365 15.355 82.535 15.525 ;
        RECT 82.365 9.915 82.535 10.085 ;
        RECT 82.825 58.875 82.995 59.045 ;
        RECT 82.825 53.435 82.995 53.605 ;
        RECT 82.825 47.995 82.995 48.165 ;
        RECT 82.825 42.555 82.995 42.725 ;
        RECT 82.825 37.115 82.995 37.285 ;
        RECT 82.825 31.675 82.995 31.845 ;
        RECT 82.825 26.235 82.995 26.405 ;
        RECT 82.825 20.795 82.995 20.965 ;
        RECT 82.825 15.355 82.995 15.525 ;
        RECT 82.825 9.915 82.995 10.085 ;
        RECT 83.285 58.875 83.455 59.045 ;
        RECT 83.285 53.435 83.455 53.605 ;
        RECT 83.285 47.995 83.455 48.165 ;
        RECT 83.285 42.555 83.455 42.725 ;
        RECT 83.285 37.115 83.455 37.285 ;
        RECT 83.285 31.675 83.455 31.845 ;
        RECT 83.285 26.235 83.455 26.405 ;
        RECT 83.285 20.795 83.455 20.965 ;
        RECT 83.285 15.355 83.455 15.525 ;
        RECT 83.285 9.915 83.455 10.085 ;
        RECT 83.745 58.875 83.915 59.045 ;
        RECT 83.745 53.435 83.915 53.605 ;
        RECT 83.745 47.995 83.915 48.165 ;
        RECT 83.745 42.555 83.915 42.725 ;
        RECT 83.745 37.115 83.915 37.285 ;
        RECT 83.745 31.675 83.915 31.845 ;
        RECT 83.745 26.235 83.915 26.405 ;
        RECT 83.745 20.795 83.915 20.965 ;
        RECT 83.745 15.355 83.915 15.525 ;
        RECT 83.745 9.915 83.915 10.085 ;
        RECT 84.205 58.875 84.375 59.045 ;
        RECT 84.205 53.435 84.375 53.605 ;
        RECT 84.205 47.995 84.375 48.165 ;
        RECT 84.205 42.555 84.375 42.725 ;
        RECT 84.205 37.115 84.375 37.285 ;
        RECT 84.205 31.675 84.375 31.845 ;
        RECT 84.205 26.235 84.375 26.405 ;
        RECT 84.205 20.795 84.375 20.965 ;
        RECT 84.205 15.355 84.375 15.525 ;
        RECT 84.205 9.915 84.375 10.085 ;
        RECT 84.665 58.875 84.835 59.045 ;
        RECT 84.665 53.435 84.835 53.605 ;
        RECT 84.665 47.995 84.835 48.165 ;
        RECT 84.665 42.555 84.835 42.725 ;
        RECT 84.665 37.115 84.835 37.285 ;
        RECT 84.665 31.675 84.835 31.845 ;
        RECT 84.665 26.235 84.835 26.405 ;
        RECT 84.665 20.795 84.835 20.965 ;
        RECT 84.665 15.355 84.835 15.525 ;
        RECT 84.665 9.915 84.835 10.085 ;
        RECT 85.125 58.875 85.295 59.045 ;
        RECT 85.125 53.435 85.295 53.605 ;
        RECT 85.125 47.995 85.295 48.165 ;
        RECT 85.125 42.555 85.295 42.725 ;
        RECT 85.125 37.115 85.295 37.285 ;
        RECT 85.125 31.675 85.295 31.845 ;
        RECT 85.125 26.235 85.295 26.405 ;
        RECT 85.125 20.795 85.295 20.965 ;
        RECT 85.125 15.355 85.295 15.525 ;
        RECT 85.125 9.915 85.295 10.085 ;
        RECT 85.585 58.875 85.755 59.045 ;
        RECT 85.585 53.435 85.755 53.605 ;
        RECT 85.585 47.995 85.755 48.165 ;
        RECT 85.585 42.555 85.755 42.725 ;
        RECT 85.585 37.115 85.755 37.285 ;
        RECT 85.585 31.675 85.755 31.845 ;
        RECT 85.585 26.235 85.755 26.405 ;
        RECT 85.585 20.795 85.755 20.965 ;
        RECT 85.585 15.355 85.755 15.525 ;
        RECT 85.585 9.915 85.755 10.085 ;
        RECT 86.045 58.875 86.215 59.045 ;
        RECT 86.045 53.435 86.215 53.605 ;
        RECT 86.045 47.995 86.215 48.165 ;
        RECT 86.045 42.555 86.215 42.725 ;
        RECT 86.045 37.115 86.215 37.285 ;
        RECT 86.045 31.675 86.215 31.845 ;
        RECT 86.045 26.235 86.215 26.405 ;
        RECT 86.045 20.795 86.215 20.965 ;
        RECT 86.045 15.355 86.215 15.525 ;
        RECT 86.045 9.915 86.215 10.085 ;
        RECT 86.505 58.875 86.675 59.045 ;
        RECT 86.505 53.435 86.675 53.605 ;
        RECT 86.505 47.995 86.675 48.165 ;
        RECT 86.505 42.555 86.675 42.725 ;
        RECT 86.505 37.115 86.675 37.285 ;
        RECT 86.505 31.675 86.675 31.845 ;
        RECT 86.505 26.235 86.675 26.405 ;
        RECT 86.505 20.795 86.675 20.965 ;
        RECT 86.505 15.355 86.675 15.525 ;
        RECT 86.505 9.915 86.675 10.085 ;
        RECT 86.965 58.875 87.135 59.045 ;
        RECT 86.965 53.435 87.135 53.605 ;
        RECT 86.965 47.995 87.135 48.165 ;
        RECT 86.965 42.555 87.135 42.725 ;
        RECT 86.965 37.115 87.135 37.285 ;
        RECT 86.965 31.675 87.135 31.845 ;
        RECT 86.965 26.235 87.135 26.405 ;
        RECT 86.965 20.795 87.135 20.965 ;
        RECT 86.965 15.355 87.135 15.525 ;
        RECT 86.965 9.915 87.135 10.085 ;
        RECT 87.425 58.875 87.595 59.045 ;
        RECT 87.425 53.435 87.595 53.605 ;
        RECT 87.425 47.995 87.595 48.165 ;
        RECT 87.425 42.555 87.595 42.725 ;
        RECT 87.425 37.115 87.595 37.285 ;
        RECT 87.425 31.675 87.595 31.845 ;
        RECT 87.425 26.235 87.595 26.405 ;
        RECT 87.425 20.795 87.595 20.965 ;
        RECT 87.425 15.355 87.595 15.525 ;
        RECT 87.425 9.915 87.595 10.085 ;
        RECT 87.885 58.875 88.055 59.045 ;
        RECT 87.885 53.435 88.055 53.605 ;
        RECT 87.885 47.995 88.055 48.165 ;
        RECT 87.885 42.555 88.055 42.725 ;
        RECT 87.885 37.115 88.055 37.285 ;
        RECT 87.885 31.675 88.055 31.845 ;
        RECT 87.885 26.235 88.055 26.405 ;
        RECT 87.885 20.795 88.055 20.965 ;
        RECT 87.885 15.355 88.055 15.525 ;
        RECT 87.885 9.915 88.055 10.085 ;
        RECT 88.345 58.875 88.515 59.045 ;
        RECT 88.345 53.435 88.515 53.605 ;
        RECT 88.345 47.995 88.515 48.165 ;
        RECT 88.345 42.555 88.515 42.725 ;
        RECT 88.345 37.115 88.515 37.285 ;
        RECT 88.345 31.675 88.515 31.845 ;
        RECT 88.345 26.235 88.515 26.405 ;
        RECT 88.345 20.795 88.515 20.965 ;
        RECT 88.345 15.355 88.515 15.525 ;
        RECT 88.345 9.915 88.515 10.085 ;
        RECT 88.805 58.875 88.975 59.045 ;
        RECT 88.805 53.435 88.975 53.605 ;
        RECT 88.805 47.995 88.975 48.165 ;
        RECT 88.805 42.555 88.975 42.725 ;
        RECT 88.805 37.115 88.975 37.285 ;
        RECT 88.805 31.675 88.975 31.845 ;
        RECT 88.805 26.235 88.975 26.405 ;
        RECT 88.805 20.795 88.975 20.965 ;
        RECT 88.805 15.355 88.975 15.525 ;
        RECT 88.805 9.915 88.975 10.085 ;
        RECT 89.265 58.875 89.435 59.045 ;
        RECT 89.265 53.435 89.435 53.605 ;
        RECT 89.265 47.995 89.435 48.165 ;
        RECT 89.265 42.555 89.435 42.725 ;
        RECT 89.265 37.115 89.435 37.285 ;
        RECT 89.265 31.675 89.435 31.845 ;
        RECT 89.265 26.235 89.435 26.405 ;
        RECT 89.265 20.795 89.435 20.965 ;
        RECT 89.265 15.355 89.435 15.525 ;
        RECT 89.265 9.915 89.435 10.085 ;
        RECT 89.725 58.875 89.895 59.045 ;
        RECT 89.725 53.435 89.895 53.605 ;
        RECT 89.725 47.995 89.895 48.165 ;
        RECT 89.725 42.555 89.895 42.725 ;
        RECT 89.725 37.115 89.895 37.285 ;
        RECT 89.725 31.675 89.895 31.845 ;
        RECT 89.725 26.235 89.895 26.405 ;
        RECT 89.725 20.795 89.895 20.965 ;
        RECT 89.725 15.355 89.895 15.525 ;
        RECT 89.725 9.915 89.895 10.085 ;
        RECT 90.185 58.875 90.355 59.045 ;
        RECT 90.185 53.435 90.355 53.605 ;
        RECT 90.185 47.995 90.355 48.165 ;
        RECT 90.185 42.555 90.355 42.725 ;
        RECT 90.185 37.115 90.355 37.285 ;
        RECT 90.185 31.675 90.355 31.845 ;
        RECT 90.185 26.235 90.355 26.405 ;
        RECT 90.185 20.795 90.355 20.965 ;
        RECT 90.185 15.355 90.355 15.525 ;
        RECT 90.185 9.915 90.355 10.085 ;
        RECT 90.645 58.875 90.815 59.045 ;
        RECT 90.645 53.435 90.815 53.605 ;
        RECT 90.645 47.995 90.815 48.165 ;
        RECT 90.645 42.555 90.815 42.725 ;
        RECT 90.645 37.115 90.815 37.285 ;
        RECT 90.645 31.675 90.815 31.845 ;
        RECT 90.645 26.235 90.815 26.405 ;
        RECT 90.645 20.795 90.815 20.965 ;
        RECT 90.645 15.355 90.815 15.525 ;
        RECT 90.645 9.915 90.815 10.085 ;
        RECT 91.105 58.875 91.275 59.045 ;
        RECT 91.105 53.435 91.275 53.605 ;
        RECT 91.105 47.995 91.275 48.165 ;
        RECT 91.105 42.555 91.275 42.725 ;
        RECT 91.105 37.115 91.275 37.285 ;
        RECT 91.105 31.675 91.275 31.845 ;
        RECT 91.105 26.235 91.275 26.405 ;
        RECT 91.105 20.795 91.275 20.965 ;
        RECT 91.105 15.355 91.275 15.525 ;
        RECT 91.105 9.915 91.275 10.085 ;
        RECT 91.565 58.875 91.735 59.045 ;
        RECT 91.565 53.435 91.735 53.605 ;
        RECT 91.565 47.995 91.735 48.165 ;
        RECT 91.565 42.555 91.735 42.725 ;
        RECT 91.565 37.115 91.735 37.285 ;
        RECT 91.565 31.675 91.735 31.845 ;
        RECT 91.565 26.235 91.735 26.405 ;
        RECT 91.565 20.795 91.735 20.965 ;
        RECT 91.565 15.355 91.735 15.525 ;
        RECT 91.565 9.915 91.735 10.085 ;
        RECT 92.025 58.875 92.195 59.045 ;
        RECT 92.025 53.435 92.195 53.605 ;
        RECT 92.025 47.995 92.195 48.165 ;
        RECT 92.025 42.555 92.195 42.725 ;
        RECT 92.025 37.115 92.195 37.285 ;
        RECT 92.025 31.675 92.195 31.845 ;
        RECT 92.025 26.235 92.195 26.405 ;
        RECT 92.025 20.795 92.195 20.965 ;
        RECT 92.025 15.355 92.195 15.525 ;
        RECT 92.025 9.915 92.195 10.085 ;
        RECT 92.485 58.875 92.655 59.045 ;
        RECT 92.485 53.435 92.655 53.605 ;
        RECT 92.485 47.995 92.655 48.165 ;
        RECT 92.485 42.555 92.655 42.725 ;
        RECT 92.485 37.115 92.655 37.285 ;
        RECT 92.485 31.675 92.655 31.845 ;
        RECT 92.485 26.235 92.655 26.405 ;
        RECT 92.485 20.795 92.655 20.965 ;
        RECT 92.485 15.355 92.655 15.525 ;
        RECT 92.485 9.915 92.655 10.085 ;
        RECT 92.945 58.875 93.115 59.045 ;
        RECT 92.945 53.435 93.115 53.605 ;
        RECT 92.945 47.995 93.115 48.165 ;
        RECT 92.945 42.555 93.115 42.725 ;
        RECT 92.945 37.115 93.115 37.285 ;
        RECT 92.945 31.675 93.115 31.845 ;
        RECT 92.945 26.235 93.115 26.405 ;
        RECT 92.945 20.795 93.115 20.965 ;
        RECT 92.945 15.355 93.115 15.525 ;
        RECT 92.945 9.915 93.115 10.085 ;
        RECT 93.405 58.875 93.575 59.045 ;
        RECT 93.405 53.435 93.575 53.605 ;
        RECT 93.405 47.995 93.575 48.165 ;
        RECT 93.405 42.555 93.575 42.725 ;
        RECT 93.405 37.115 93.575 37.285 ;
        RECT 93.405 31.675 93.575 31.845 ;
        RECT 93.405 26.235 93.575 26.405 ;
        RECT 93.405 20.795 93.575 20.965 ;
        RECT 93.405 15.355 93.575 15.525 ;
        RECT 93.405 9.915 93.575 10.085 ;
        RECT 93.865 58.875 94.035 59.045 ;
        RECT 93.865 53.435 94.035 53.605 ;
        RECT 93.865 47.995 94.035 48.165 ;
        RECT 93.865 42.555 94.035 42.725 ;
        RECT 93.865 37.115 94.035 37.285 ;
        RECT 93.865 31.675 94.035 31.845 ;
        RECT 93.865 26.235 94.035 26.405 ;
        RECT 93.865 20.795 94.035 20.965 ;
        RECT 93.865 15.355 94.035 15.525 ;
        RECT 93.865 9.915 94.035 10.085 ;
        RECT 94.325 58.875 94.495 59.045 ;
        RECT 94.325 53.435 94.495 53.605 ;
        RECT 94.325 47.995 94.495 48.165 ;
        RECT 94.325 42.555 94.495 42.725 ;
        RECT 94.325 37.115 94.495 37.285 ;
        RECT 94.325 31.675 94.495 31.845 ;
        RECT 94.325 26.235 94.495 26.405 ;
        RECT 94.325 20.795 94.495 20.965 ;
        RECT 94.325 15.355 94.495 15.525 ;
        RECT 94.325 9.915 94.495 10.085 ;
        RECT 94.785 58.875 94.955 59.045 ;
        RECT 94.785 53.435 94.955 53.605 ;
        RECT 94.785 47.995 94.955 48.165 ;
        RECT 94.785 42.555 94.955 42.725 ;
        RECT 94.785 37.115 94.955 37.285 ;
        RECT 94.785 31.675 94.955 31.845 ;
        RECT 94.785 26.235 94.955 26.405 ;
        RECT 94.785 20.795 94.955 20.965 ;
        RECT 94.785 15.355 94.955 15.525 ;
        RECT 94.785 9.915 94.955 10.085 ;
        RECT 95.245 58.875 95.415 59.045 ;
        RECT 95.245 53.435 95.415 53.605 ;
        RECT 95.245 47.995 95.415 48.165 ;
        RECT 95.245 42.555 95.415 42.725 ;
        RECT 95.245 37.115 95.415 37.285 ;
        RECT 95.245 31.675 95.415 31.845 ;
        RECT 95.245 26.235 95.415 26.405 ;
        RECT 95.245 20.795 95.415 20.965 ;
        RECT 95.245 15.355 95.415 15.525 ;
        RECT 95.245 9.915 95.415 10.085 ;
        RECT 95.705 58.875 95.875 59.045 ;
        RECT 95.705 53.435 95.875 53.605 ;
        RECT 95.705 47.995 95.875 48.165 ;
        RECT 95.705 42.555 95.875 42.725 ;
        RECT 95.705 37.115 95.875 37.285 ;
        RECT 95.705 31.675 95.875 31.845 ;
        RECT 95.705 26.235 95.875 26.405 ;
        RECT 95.705 20.795 95.875 20.965 ;
        RECT 95.705 15.355 95.875 15.525 ;
        RECT 95.705 9.915 95.875 10.085 ;
        RECT 96.165 58.875 96.335 59.045 ;
        RECT 96.165 53.435 96.335 53.605 ;
        RECT 96.165 47.995 96.335 48.165 ;
        RECT 96.165 42.555 96.335 42.725 ;
        RECT 96.165 37.115 96.335 37.285 ;
        RECT 96.165 31.675 96.335 31.845 ;
        RECT 96.165 26.235 96.335 26.405 ;
        RECT 96.165 20.795 96.335 20.965 ;
        RECT 96.165 15.355 96.335 15.525 ;
        RECT 96.165 9.915 96.335 10.085 ;
        RECT 96.625 58.875 96.795 59.045 ;
        RECT 96.625 53.435 96.795 53.605 ;
        RECT 96.625 47.995 96.795 48.165 ;
        RECT 96.625 42.555 96.795 42.725 ;
        RECT 96.625 37.115 96.795 37.285 ;
        RECT 96.625 31.675 96.795 31.845 ;
        RECT 96.625 26.235 96.795 26.405 ;
        RECT 96.625 20.795 96.795 20.965 ;
        RECT 96.625 15.355 96.795 15.525 ;
        RECT 96.625 9.915 96.795 10.085 ;
        RECT 97.085 58.875 97.255 59.045 ;
        RECT 97.085 53.435 97.255 53.605 ;
        RECT 97.085 47.995 97.255 48.165 ;
        RECT 97.085 42.555 97.255 42.725 ;
        RECT 97.085 37.115 97.255 37.285 ;
        RECT 97.085 31.675 97.255 31.845 ;
        RECT 97.085 26.235 97.255 26.405 ;
        RECT 97.085 20.795 97.255 20.965 ;
        RECT 97.085 15.355 97.255 15.525 ;
        RECT 97.085 9.915 97.255 10.085 ;
        RECT 97.545 58.875 97.715 59.045 ;
        RECT 97.545 53.435 97.715 53.605 ;
        RECT 97.545 47.995 97.715 48.165 ;
        RECT 97.545 42.555 97.715 42.725 ;
        RECT 97.545 37.115 97.715 37.285 ;
        RECT 97.545 31.675 97.715 31.845 ;
        RECT 97.545 26.235 97.715 26.405 ;
        RECT 97.545 20.795 97.715 20.965 ;
        RECT 97.545 15.355 97.715 15.525 ;
        RECT 97.545 9.915 97.715 10.085 ;
        RECT 98.005 58.875 98.175 59.045 ;
        RECT 98.005 53.435 98.175 53.605 ;
        RECT 98.005 47.995 98.175 48.165 ;
        RECT 98.005 42.555 98.175 42.725 ;
        RECT 98.005 37.115 98.175 37.285 ;
        RECT 98.005 31.675 98.175 31.845 ;
        RECT 98.005 26.235 98.175 26.405 ;
        RECT 98.005 20.795 98.175 20.965 ;
        RECT 98.005 15.355 98.175 15.525 ;
        RECT 98.005 9.915 98.175 10.085 ;
        RECT 98.465 58.875 98.635 59.045 ;
        RECT 98.465 53.435 98.635 53.605 ;
        RECT 98.465 47.995 98.635 48.165 ;
        RECT 98.465 42.555 98.635 42.725 ;
        RECT 98.465 37.115 98.635 37.285 ;
        RECT 98.465 31.675 98.635 31.845 ;
        RECT 98.465 26.235 98.635 26.405 ;
        RECT 98.465 20.795 98.635 20.965 ;
        RECT 98.465 15.355 98.635 15.525 ;
        RECT 98.465 9.915 98.635 10.085 ;
        RECT 98.925 58.875 99.095 59.045 ;
        RECT 98.925 53.435 99.095 53.605 ;
        RECT 98.925 47.995 99.095 48.165 ;
        RECT 98.925 42.555 99.095 42.725 ;
        RECT 98.925 37.115 99.095 37.285 ;
        RECT 98.925 31.675 99.095 31.845 ;
        RECT 98.925 26.235 99.095 26.405 ;
        RECT 98.925 20.795 99.095 20.965 ;
        RECT 98.925 15.355 99.095 15.525 ;
        RECT 98.925 9.915 99.095 10.085 ;
        RECT 99.385 58.875 99.555 59.045 ;
        RECT 99.385 53.435 99.555 53.605 ;
        RECT 99.385 47.995 99.555 48.165 ;
        RECT 99.385 42.555 99.555 42.725 ;
        RECT 99.385 37.115 99.555 37.285 ;
        RECT 99.385 31.675 99.555 31.845 ;
        RECT 99.385 26.235 99.555 26.405 ;
        RECT 99.385 20.795 99.555 20.965 ;
        RECT 99.385 15.355 99.555 15.525 ;
        RECT 99.385 9.915 99.555 10.085 ;
        RECT 99.845 58.875 100.015 59.045 ;
        RECT 99.845 53.435 100.015 53.605 ;
        RECT 99.845 47.995 100.015 48.165 ;
        RECT 99.845 42.555 100.015 42.725 ;
        RECT 99.845 37.115 100.015 37.285 ;
        RECT 99.845 31.675 100.015 31.845 ;
        RECT 99.845 26.235 100.015 26.405 ;
        RECT 99.845 20.795 100.015 20.965 ;
        RECT 99.845 15.355 100.015 15.525 ;
        RECT 99.845 9.915 100.015 10.085 ;
        RECT 100.305 58.875 100.475 59.045 ;
        RECT 100.305 53.435 100.475 53.605 ;
        RECT 100.305 47.995 100.475 48.165 ;
        RECT 100.305 42.555 100.475 42.725 ;
        RECT 100.305 37.115 100.475 37.285 ;
        RECT 100.305 31.675 100.475 31.845 ;
        RECT 100.305 26.235 100.475 26.405 ;
        RECT 100.305 20.795 100.475 20.965 ;
        RECT 100.305 15.355 100.475 15.525 ;
        RECT 100.305 9.915 100.475 10.085 ;
        RECT 100.765 58.875 100.935 59.045 ;
        RECT 100.765 53.435 100.935 53.605 ;
        RECT 100.765 47.995 100.935 48.165 ;
        RECT 100.765 42.555 100.935 42.725 ;
        RECT 100.765 37.115 100.935 37.285 ;
        RECT 100.765 31.675 100.935 31.845 ;
        RECT 100.765 26.235 100.935 26.405 ;
        RECT 100.765 20.795 100.935 20.965 ;
        RECT 100.765 15.355 100.935 15.525 ;
        RECT 100.765 9.915 100.935 10.085 ;
        RECT 101.225 58.875 101.395 59.045 ;
        RECT 101.225 53.435 101.395 53.605 ;
        RECT 101.225 47.995 101.395 48.165 ;
        RECT 101.225 42.555 101.395 42.725 ;
        RECT 101.225 37.115 101.395 37.285 ;
        RECT 101.225 31.675 101.395 31.845 ;
        RECT 101.225 26.235 101.395 26.405 ;
        RECT 101.225 20.795 101.395 20.965 ;
        RECT 101.225 15.355 101.395 15.525 ;
        RECT 101.225 9.915 101.395 10.085 ;
        RECT 101.685 58.875 101.855 59.045 ;
        RECT 101.685 53.435 101.855 53.605 ;
        RECT 101.685 47.995 101.855 48.165 ;
        RECT 101.685 42.555 101.855 42.725 ;
        RECT 101.685 37.115 101.855 37.285 ;
        RECT 101.685 31.675 101.855 31.845 ;
        RECT 101.685 26.235 101.855 26.405 ;
        RECT 101.685 20.795 101.855 20.965 ;
        RECT 101.685 15.355 101.855 15.525 ;
        RECT 101.685 9.915 101.855 10.085 ;
        RECT 10.145 58.875 10.315 59.045 ;
        RECT 10.145 53.435 10.315 53.605 ;
        RECT 10.145 47.995 10.315 48.165 ;
        RECT 10.145 42.555 10.315 42.725 ;
        RECT 10.145 37.115 10.315 37.285 ;
        RECT 10.145 31.675 10.315 31.845 ;
        RECT 10.145 26.235 10.315 26.405 ;
        RECT 10.145 20.795 10.315 20.965 ;
        RECT 10.145 15.355 10.315 15.525 ;
        RECT 10.145 9.915 10.315 10.085 ;
        RECT 10.605 58.875 10.775 59.045 ;
        RECT 10.605 53.435 10.775 53.605 ;
        RECT 10.605 47.995 10.775 48.165 ;
        RECT 10.605 42.555 10.775 42.725 ;
        RECT 10.605 37.115 10.775 37.285 ;
        RECT 10.605 31.675 10.775 31.845 ;
        RECT 10.605 26.235 10.775 26.405 ;
        RECT 10.605 20.795 10.775 20.965 ;
        RECT 10.605 15.355 10.775 15.525 ;
        RECT 10.605 9.915 10.775 10.085 ;
        RECT 11.065 58.875 11.235 59.045 ;
        RECT 11.065 53.435 11.235 53.605 ;
        RECT 11.065 47.995 11.235 48.165 ;
        RECT 11.065 42.555 11.235 42.725 ;
        RECT 11.065 37.115 11.235 37.285 ;
        RECT 11.065 31.675 11.235 31.845 ;
        RECT 11.065 26.235 11.235 26.405 ;
        RECT 11.065 20.795 11.235 20.965 ;
        RECT 11.065 15.355 11.235 15.525 ;
        RECT 11.065 9.915 11.235 10.085 ;
        RECT 11.525 58.875 11.695 59.045 ;
        RECT 11.525 53.435 11.695 53.605 ;
        RECT 11.525 47.995 11.695 48.165 ;
        RECT 11.525 42.555 11.695 42.725 ;
        RECT 11.525 37.115 11.695 37.285 ;
        RECT 11.525 31.675 11.695 31.845 ;
        RECT 11.525 26.235 11.695 26.405 ;
        RECT 11.525 20.795 11.695 20.965 ;
        RECT 11.525 15.355 11.695 15.525 ;
        RECT 11.525 9.915 11.695 10.085 ;
        RECT 11.985 58.875 12.155 59.045 ;
        RECT 11.985 53.435 12.155 53.605 ;
        RECT 11.985 47.995 12.155 48.165 ;
        RECT 11.985 42.555 12.155 42.725 ;
        RECT 11.985 37.115 12.155 37.285 ;
        RECT 11.985 31.675 12.155 31.845 ;
        RECT 11.985 26.235 12.155 26.405 ;
        RECT 11.985 20.795 12.155 20.965 ;
        RECT 11.985 15.355 12.155 15.525 ;
        RECT 11.985 9.915 12.155 10.085 ;
        RECT 12.445 58.875 12.615 59.045 ;
        RECT 12.445 53.435 12.615 53.605 ;
        RECT 12.445 47.995 12.615 48.165 ;
        RECT 12.445 42.555 12.615 42.725 ;
        RECT 12.445 37.115 12.615 37.285 ;
        RECT 12.445 31.675 12.615 31.845 ;
        RECT 12.445 26.235 12.615 26.405 ;
        RECT 12.445 20.795 12.615 20.965 ;
        RECT 12.445 15.355 12.615 15.525 ;
        RECT 12.445 9.915 12.615 10.085 ;
        RECT 12.905 58.875 13.075 59.045 ;
        RECT 12.905 53.435 13.075 53.605 ;
        RECT 12.905 47.995 13.075 48.165 ;
        RECT 12.905 42.555 13.075 42.725 ;
        RECT 12.905 37.115 13.075 37.285 ;
        RECT 12.905 31.675 13.075 31.845 ;
        RECT 12.905 26.235 13.075 26.405 ;
        RECT 12.905 20.795 13.075 20.965 ;
        RECT 12.905 15.355 13.075 15.525 ;
        RECT 12.905 9.915 13.075 10.085 ;
        RECT 13.365 58.875 13.535 59.045 ;
        RECT 13.365 53.435 13.535 53.605 ;
        RECT 13.365 47.995 13.535 48.165 ;
        RECT 13.365 42.555 13.535 42.725 ;
        RECT 13.365 37.115 13.535 37.285 ;
        RECT 13.365 31.675 13.535 31.845 ;
        RECT 13.365 26.235 13.535 26.405 ;
        RECT 13.365 20.795 13.535 20.965 ;
        RECT 13.365 15.355 13.535 15.525 ;
        RECT 13.365 9.915 13.535 10.085 ;
        RECT 13.825 58.875 13.995 59.045 ;
        RECT 13.825 53.435 13.995 53.605 ;
        RECT 13.825 47.995 13.995 48.165 ;
        RECT 13.825 42.555 13.995 42.725 ;
        RECT 13.825 37.115 13.995 37.285 ;
        RECT 13.825 31.675 13.995 31.845 ;
        RECT 13.825 26.235 13.995 26.405 ;
        RECT 13.825 20.795 13.995 20.965 ;
        RECT 13.825 15.355 13.995 15.525 ;
        RECT 13.825 9.915 13.995 10.085 ;
        RECT 14.285 58.875 14.455 59.045 ;
        RECT 14.285 53.435 14.455 53.605 ;
        RECT 14.285 47.995 14.455 48.165 ;
        RECT 14.285 42.555 14.455 42.725 ;
        RECT 14.285 37.115 14.455 37.285 ;
        RECT 14.285 31.675 14.455 31.845 ;
        RECT 14.285 26.235 14.455 26.405 ;
        RECT 14.285 20.795 14.455 20.965 ;
        RECT 14.285 15.355 14.455 15.525 ;
        RECT 14.285 9.915 14.455 10.085 ;
        RECT 14.745 58.875 14.915 59.045 ;
        RECT 14.745 53.435 14.915 53.605 ;
        RECT 14.745 47.995 14.915 48.165 ;
        RECT 14.745 42.555 14.915 42.725 ;
        RECT 14.745 37.115 14.915 37.285 ;
        RECT 14.745 31.675 14.915 31.845 ;
        RECT 14.745 26.235 14.915 26.405 ;
        RECT 14.745 20.795 14.915 20.965 ;
        RECT 14.745 15.355 14.915 15.525 ;
        RECT 14.745 9.915 14.915 10.085 ;
        RECT 15.205 58.875 15.375 59.045 ;
        RECT 15.205 53.435 15.375 53.605 ;
        RECT 15.205 47.995 15.375 48.165 ;
        RECT 15.205 42.555 15.375 42.725 ;
        RECT 15.205 37.115 15.375 37.285 ;
        RECT 15.205 31.675 15.375 31.845 ;
        RECT 15.205 26.235 15.375 26.405 ;
        RECT 15.205 20.795 15.375 20.965 ;
        RECT 15.205 15.355 15.375 15.525 ;
        RECT 15.205 9.915 15.375 10.085 ;
        RECT 15.665 58.875 15.835 59.045 ;
        RECT 15.665 53.435 15.835 53.605 ;
        RECT 15.665 47.995 15.835 48.165 ;
        RECT 15.665 42.555 15.835 42.725 ;
        RECT 15.665 37.115 15.835 37.285 ;
        RECT 15.665 31.675 15.835 31.845 ;
        RECT 15.665 26.235 15.835 26.405 ;
        RECT 15.665 20.795 15.835 20.965 ;
        RECT 15.665 15.355 15.835 15.525 ;
        RECT 15.665 9.915 15.835 10.085 ;
        RECT 16.125 58.875 16.295 59.045 ;
        RECT 16.125 53.435 16.295 53.605 ;
        RECT 16.125 47.995 16.295 48.165 ;
        RECT 16.125 42.555 16.295 42.725 ;
        RECT 16.125 37.115 16.295 37.285 ;
        RECT 16.125 31.675 16.295 31.845 ;
        RECT 16.125 26.235 16.295 26.405 ;
        RECT 16.125 20.795 16.295 20.965 ;
        RECT 16.125 15.355 16.295 15.525 ;
        RECT 16.125 9.915 16.295 10.085 ;
        RECT 16.585 58.875 16.755 59.045 ;
        RECT 16.585 53.435 16.755 53.605 ;
        RECT 16.585 47.995 16.755 48.165 ;
        RECT 16.585 42.555 16.755 42.725 ;
        RECT 16.585 37.115 16.755 37.285 ;
        RECT 16.585 31.675 16.755 31.845 ;
        RECT 16.585 26.235 16.755 26.405 ;
        RECT 16.585 20.795 16.755 20.965 ;
        RECT 16.585 15.355 16.755 15.525 ;
        RECT 16.585 9.915 16.755 10.085 ;
        RECT 17.045 58.875 17.215 59.045 ;
        RECT 17.045 53.435 17.215 53.605 ;
        RECT 17.045 47.995 17.215 48.165 ;
        RECT 17.045 42.555 17.215 42.725 ;
        RECT 17.045 37.115 17.215 37.285 ;
        RECT 17.045 31.675 17.215 31.845 ;
        RECT 17.045 26.235 17.215 26.405 ;
        RECT 17.045 20.795 17.215 20.965 ;
        RECT 17.045 15.355 17.215 15.525 ;
        RECT 17.045 9.915 17.215 10.085 ;
        RECT 17.505 58.875 17.675 59.045 ;
        RECT 17.505 53.435 17.675 53.605 ;
        RECT 17.505 47.995 17.675 48.165 ;
        RECT 17.505 42.555 17.675 42.725 ;
        RECT 17.505 37.115 17.675 37.285 ;
        RECT 17.505 31.675 17.675 31.845 ;
        RECT 17.505 26.235 17.675 26.405 ;
        RECT 17.505 20.795 17.675 20.965 ;
        RECT 17.505 15.355 17.675 15.525 ;
        RECT 17.505 9.915 17.675 10.085 ;
        RECT 17.965 58.875 18.135 59.045 ;
        RECT 17.965 53.435 18.135 53.605 ;
        RECT 17.965 47.995 18.135 48.165 ;
        RECT 17.965 42.555 18.135 42.725 ;
        RECT 17.965 37.115 18.135 37.285 ;
        RECT 17.965 31.675 18.135 31.845 ;
        RECT 17.965 26.235 18.135 26.405 ;
        RECT 17.965 20.795 18.135 20.965 ;
        RECT 17.965 15.355 18.135 15.525 ;
        RECT 17.965 9.915 18.135 10.085 ;
        RECT 18.425 58.875 18.595 59.045 ;
        RECT 18.425 53.435 18.595 53.605 ;
        RECT 18.425 47.995 18.595 48.165 ;
        RECT 18.425 42.555 18.595 42.725 ;
        RECT 18.425 37.115 18.595 37.285 ;
        RECT 18.425 31.675 18.595 31.845 ;
        RECT 18.425 26.235 18.595 26.405 ;
        RECT 18.425 20.795 18.595 20.965 ;
        RECT 18.425 15.355 18.595 15.525 ;
        RECT 18.425 9.915 18.595 10.085 ;
        RECT 18.885 58.875 19.055 59.045 ;
        RECT 18.885 53.435 19.055 53.605 ;
        RECT 18.885 47.995 19.055 48.165 ;
        RECT 18.885 42.555 19.055 42.725 ;
        RECT 18.885 37.115 19.055 37.285 ;
        RECT 18.885 31.675 19.055 31.845 ;
        RECT 18.885 26.235 19.055 26.405 ;
        RECT 18.885 20.795 19.055 20.965 ;
        RECT 18.885 15.355 19.055 15.525 ;
        RECT 18.885 9.915 19.055 10.085 ;
        RECT 19.345 58.875 19.515 59.045 ;
        RECT 19.345 53.435 19.515 53.605 ;
        RECT 19.345 47.995 19.515 48.165 ;
        RECT 19.345 42.555 19.515 42.725 ;
        RECT 19.345 37.115 19.515 37.285 ;
        RECT 19.345 31.675 19.515 31.845 ;
        RECT 19.345 26.235 19.515 26.405 ;
        RECT 19.345 20.795 19.515 20.965 ;
        RECT 19.345 15.355 19.515 15.525 ;
        RECT 19.345 9.915 19.515 10.085 ;
        RECT 19.805 58.875 19.975 59.045 ;
        RECT 19.805 53.435 19.975 53.605 ;
        RECT 19.805 47.995 19.975 48.165 ;
        RECT 19.805 42.555 19.975 42.725 ;
        RECT 19.805 37.115 19.975 37.285 ;
        RECT 19.805 31.675 19.975 31.845 ;
        RECT 19.805 26.235 19.975 26.405 ;
        RECT 19.805 20.795 19.975 20.965 ;
        RECT 19.805 15.355 19.975 15.525 ;
        RECT 19.805 9.915 19.975 10.085 ;
        RECT 20.265 58.875 20.435 59.045 ;
        RECT 20.265 53.435 20.435 53.605 ;
        RECT 20.265 47.995 20.435 48.165 ;
        RECT 20.265 42.555 20.435 42.725 ;
        RECT 20.265 37.115 20.435 37.285 ;
        RECT 20.265 31.675 20.435 31.845 ;
        RECT 20.265 26.235 20.435 26.405 ;
        RECT 20.265 20.795 20.435 20.965 ;
        RECT 20.265 15.355 20.435 15.525 ;
        RECT 20.265 9.915 20.435 10.085 ;
        RECT 20.725 58.875 20.895 59.045 ;
        RECT 20.725 53.435 20.895 53.605 ;
        RECT 20.725 47.995 20.895 48.165 ;
        RECT 20.725 42.555 20.895 42.725 ;
        RECT 20.725 37.115 20.895 37.285 ;
        RECT 20.725 31.675 20.895 31.845 ;
        RECT 20.725 26.235 20.895 26.405 ;
        RECT 20.725 20.795 20.895 20.965 ;
        RECT 20.725 15.355 20.895 15.525 ;
        RECT 20.725 9.915 20.895 10.085 ;
        RECT 21.185 58.875 21.355 59.045 ;
        RECT 21.185 53.435 21.355 53.605 ;
        RECT 21.185 47.995 21.355 48.165 ;
        RECT 21.185 42.555 21.355 42.725 ;
        RECT 21.185 37.115 21.355 37.285 ;
        RECT 21.185 31.675 21.355 31.845 ;
        RECT 21.185 26.235 21.355 26.405 ;
        RECT 21.185 20.795 21.355 20.965 ;
        RECT 21.185 15.355 21.355 15.525 ;
        RECT 21.185 9.915 21.355 10.085 ;
        RECT 21.645 58.875 21.815 59.045 ;
        RECT 21.645 53.435 21.815 53.605 ;
        RECT 21.645 47.995 21.815 48.165 ;
        RECT 21.645 42.555 21.815 42.725 ;
        RECT 21.645 37.115 21.815 37.285 ;
        RECT 21.645 31.675 21.815 31.845 ;
        RECT 21.645 26.235 21.815 26.405 ;
        RECT 21.645 20.795 21.815 20.965 ;
        RECT 21.645 15.355 21.815 15.525 ;
        RECT 21.645 9.915 21.815 10.085 ;
        RECT 22.105 58.875 22.275 59.045 ;
        RECT 22.105 53.435 22.275 53.605 ;
        RECT 22.105 47.995 22.275 48.165 ;
        RECT 22.105 42.555 22.275 42.725 ;
        RECT 22.105 37.115 22.275 37.285 ;
        RECT 22.105 31.675 22.275 31.845 ;
        RECT 22.105 26.235 22.275 26.405 ;
        RECT 22.105 20.795 22.275 20.965 ;
        RECT 22.105 15.355 22.275 15.525 ;
        RECT 22.105 9.915 22.275 10.085 ;
        RECT 22.565 58.875 22.735 59.045 ;
        RECT 22.565 53.435 22.735 53.605 ;
        RECT 22.565 47.995 22.735 48.165 ;
        RECT 22.565 42.555 22.735 42.725 ;
        RECT 22.565 37.115 22.735 37.285 ;
        RECT 22.565 31.675 22.735 31.845 ;
        RECT 22.565 26.235 22.735 26.405 ;
        RECT 22.565 20.795 22.735 20.965 ;
        RECT 22.565 15.355 22.735 15.525 ;
        RECT 22.565 9.915 22.735 10.085 ;
        RECT 23.025 58.875 23.195 59.045 ;
        RECT 23.025 53.435 23.195 53.605 ;
        RECT 23.025 47.995 23.195 48.165 ;
        RECT 23.025 42.555 23.195 42.725 ;
        RECT 23.025 37.115 23.195 37.285 ;
        RECT 23.025 31.675 23.195 31.845 ;
        RECT 23.025 26.235 23.195 26.405 ;
        RECT 23.025 20.795 23.195 20.965 ;
        RECT 23.025 15.355 23.195 15.525 ;
        RECT 23.025 9.915 23.195 10.085 ;
        RECT 23.485 58.875 23.655 59.045 ;
        RECT 23.485 53.435 23.655 53.605 ;
        RECT 23.485 47.995 23.655 48.165 ;
        RECT 23.485 42.555 23.655 42.725 ;
        RECT 23.485 37.115 23.655 37.285 ;
        RECT 23.485 31.675 23.655 31.845 ;
        RECT 23.485 26.235 23.655 26.405 ;
        RECT 23.485 20.795 23.655 20.965 ;
        RECT 23.485 15.355 23.655 15.525 ;
        RECT 23.485 9.915 23.655 10.085 ;
        RECT 23.945 58.875 24.115 59.045 ;
        RECT 23.945 53.435 24.115 53.605 ;
        RECT 23.945 47.995 24.115 48.165 ;
        RECT 23.945 42.555 24.115 42.725 ;
        RECT 23.945 37.115 24.115 37.285 ;
        RECT 23.945 31.675 24.115 31.845 ;
        RECT 23.945 26.235 24.115 26.405 ;
        RECT 23.945 20.795 24.115 20.965 ;
        RECT 23.945 15.355 24.115 15.525 ;
        RECT 23.945 9.915 24.115 10.085 ;
        RECT 24.405 58.875 24.575 59.045 ;
        RECT 24.405 53.435 24.575 53.605 ;
        RECT 24.405 47.995 24.575 48.165 ;
        RECT 24.405 42.555 24.575 42.725 ;
        RECT 24.405 37.115 24.575 37.285 ;
        RECT 24.405 31.675 24.575 31.845 ;
        RECT 24.405 26.235 24.575 26.405 ;
        RECT 24.405 20.795 24.575 20.965 ;
        RECT 24.405 15.355 24.575 15.525 ;
        RECT 24.405 9.915 24.575 10.085 ;
        RECT 24.865 58.875 25.035 59.045 ;
        RECT 24.865 53.435 25.035 53.605 ;
        RECT 24.865 47.995 25.035 48.165 ;
        RECT 24.865 42.555 25.035 42.725 ;
        RECT 24.865 37.115 25.035 37.285 ;
        RECT 24.865 31.675 25.035 31.845 ;
        RECT 24.865 26.235 25.035 26.405 ;
        RECT 24.865 20.795 25.035 20.965 ;
        RECT 24.865 15.355 25.035 15.525 ;
        RECT 24.865 9.915 25.035 10.085 ;
        RECT 25.325 58.875 25.495 59.045 ;
        RECT 25.325 53.435 25.495 53.605 ;
        RECT 25.325 47.995 25.495 48.165 ;
        RECT 25.325 42.555 25.495 42.725 ;
        RECT 25.325 37.115 25.495 37.285 ;
        RECT 25.325 31.675 25.495 31.845 ;
        RECT 25.325 26.235 25.495 26.405 ;
        RECT 25.325 20.795 25.495 20.965 ;
        RECT 25.325 15.355 25.495 15.525 ;
        RECT 25.325 9.915 25.495 10.085 ;
        RECT 25.785 58.875 25.955 59.045 ;
        RECT 25.785 53.435 25.955 53.605 ;
        RECT 25.785 47.995 25.955 48.165 ;
        RECT 25.785 42.555 25.955 42.725 ;
        RECT 25.785 37.115 25.955 37.285 ;
        RECT 25.785 31.675 25.955 31.845 ;
        RECT 25.785 26.235 25.955 26.405 ;
        RECT 25.785 20.795 25.955 20.965 ;
        RECT 25.785 15.355 25.955 15.525 ;
        RECT 25.785 9.915 25.955 10.085 ;
        RECT 26.245 58.875 26.415 59.045 ;
        RECT 26.245 53.435 26.415 53.605 ;
        RECT 26.245 47.995 26.415 48.165 ;
        RECT 26.245 42.555 26.415 42.725 ;
        RECT 26.245 37.115 26.415 37.285 ;
        RECT 26.245 31.675 26.415 31.845 ;
        RECT 26.245 26.235 26.415 26.405 ;
        RECT 26.245 20.795 26.415 20.965 ;
        RECT 26.245 15.355 26.415 15.525 ;
        RECT 26.245 9.915 26.415 10.085 ;
        RECT 26.705 58.875 26.875 59.045 ;
        RECT 26.705 53.435 26.875 53.605 ;
        RECT 26.705 47.995 26.875 48.165 ;
        RECT 26.705 42.555 26.875 42.725 ;
        RECT 26.705 37.115 26.875 37.285 ;
        RECT 26.705 31.675 26.875 31.845 ;
        RECT 26.705 26.235 26.875 26.405 ;
        RECT 26.705 20.795 26.875 20.965 ;
        RECT 26.705 15.355 26.875 15.525 ;
        RECT 26.705 9.915 26.875 10.085 ;
        RECT 27.165 58.875 27.335 59.045 ;
        RECT 27.165 53.435 27.335 53.605 ;
        RECT 27.165 47.995 27.335 48.165 ;
        RECT 27.165 42.555 27.335 42.725 ;
        RECT 27.165 37.115 27.335 37.285 ;
        RECT 27.165 31.675 27.335 31.845 ;
        RECT 27.165 26.235 27.335 26.405 ;
        RECT 27.165 20.795 27.335 20.965 ;
        RECT 27.165 15.355 27.335 15.525 ;
        RECT 27.165 9.915 27.335 10.085 ;
        RECT 27.625 58.875 27.795 59.045 ;
        RECT 27.625 53.435 27.795 53.605 ;
        RECT 27.625 47.995 27.795 48.165 ;
        RECT 27.625 42.555 27.795 42.725 ;
        RECT 27.625 37.115 27.795 37.285 ;
        RECT 27.625 31.675 27.795 31.845 ;
        RECT 27.625 26.235 27.795 26.405 ;
        RECT 27.625 20.795 27.795 20.965 ;
        RECT 27.625 15.355 27.795 15.525 ;
        RECT 27.625 9.915 27.795 10.085 ;
        RECT 28.085 58.875 28.255 59.045 ;
        RECT 28.085 53.435 28.255 53.605 ;
        RECT 28.085 47.995 28.255 48.165 ;
        RECT 28.085 42.555 28.255 42.725 ;
        RECT 28.085 37.115 28.255 37.285 ;
        RECT 28.085 31.675 28.255 31.845 ;
        RECT 28.085 26.235 28.255 26.405 ;
        RECT 28.085 20.795 28.255 20.965 ;
        RECT 28.085 15.355 28.255 15.525 ;
        RECT 28.085 9.915 28.255 10.085 ;
        RECT 28.545 58.875 28.715 59.045 ;
        RECT 28.545 53.435 28.715 53.605 ;
        RECT 28.545 47.995 28.715 48.165 ;
        RECT 28.545 42.555 28.715 42.725 ;
        RECT 28.545 37.115 28.715 37.285 ;
        RECT 28.545 31.675 28.715 31.845 ;
        RECT 28.545 26.235 28.715 26.405 ;
        RECT 28.545 20.795 28.715 20.965 ;
        RECT 28.545 15.355 28.715 15.525 ;
        RECT 28.545 9.915 28.715 10.085 ;
        RECT 29.005 58.875 29.175 59.045 ;
        RECT 29.005 53.435 29.175 53.605 ;
        RECT 29.005 47.995 29.175 48.165 ;
        RECT 29.005 42.555 29.175 42.725 ;
        RECT 29.005 37.115 29.175 37.285 ;
        RECT 29.005 31.675 29.175 31.845 ;
        RECT 29.005 26.235 29.175 26.405 ;
        RECT 29.005 20.795 29.175 20.965 ;
        RECT 29.005 15.355 29.175 15.525 ;
        RECT 29.005 9.915 29.175 10.085 ;
        RECT 29.465 58.875 29.635 59.045 ;
        RECT 29.465 53.435 29.635 53.605 ;
        RECT 29.465 47.995 29.635 48.165 ;
        RECT 29.465 42.555 29.635 42.725 ;
        RECT 29.465 37.115 29.635 37.285 ;
        RECT 29.465 31.675 29.635 31.845 ;
        RECT 29.465 26.235 29.635 26.405 ;
        RECT 29.465 20.795 29.635 20.965 ;
        RECT 29.465 15.355 29.635 15.525 ;
        RECT 29.465 9.915 29.635 10.085 ;
        RECT 29.925 58.875 30.095 59.045 ;
        RECT 29.925 53.435 30.095 53.605 ;
        RECT 29.925 47.995 30.095 48.165 ;
        RECT 29.925 42.555 30.095 42.725 ;
        RECT 29.925 37.115 30.095 37.285 ;
        RECT 29.925 31.675 30.095 31.845 ;
        RECT 29.925 26.235 30.095 26.405 ;
        RECT 29.925 20.795 30.095 20.965 ;
        RECT 29.925 15.355 30.095 15.525 ;
        RECT 29.925 9.915 30.095 10.085 ;
        RECT 30.385 58.875 30.555 59.045 ;
        RECT 30.385 53.435 30.555 53.605 ;
        RECT 30.385 47.995 30.555 48.165 ;
        RECT 30.385 42.555 30.555 42.725 ;
        RECT 30.385 37.115 30.555 37.285 ;
        RECT 30.385 31.675 30.555 31.845 ;
        RECT 30.385 26.235 30.555 26.405 ;
        RECT 30.385 20.795 30.555 20.965 ;
        RECT 30.385 15.355 30.555 15.525 ;
        RECT 30.385 9.915 30.555 10.085 ;
        RECT 30.845 58.875 31.015 59.045 ;
        RECT 30.845 53.435 31.015 53.605 ;
        RECT 30.845 47.995 31.015 48.165 ;
        RECT 30.845 42.555 31.015 42.725 ;
        RECT 30.845 37.115 31.015 37.285 ;
        RECT 30.845 31.675 31.015 31.845 ;
        RECT 30.845 26.235 31.015 26.405 ;
        RECT 30.845 20.795 31.015 20.965 ;
        RECT 30.845 15.355 31.015 15.525 ;
        RECT 30.845 9.915 31.015 10.085 ;
        RECT 31.305 58.875 31.475 59.045 ;
        RECT 31.305 53.435 31.475 53.605 ;
        RECT 31.305 47.995 31.475 48.165 ;
        RECT 31.305 42.555 31.475 42.725 ;
        RECT 31.305 37.115 31.475 37.285 ;
        RECT 31.305 31.675 31.475 31.845 ;
        RECT 31.305 26.235 31.475 26.405 ;
        RECT 31.305 20.795 31.475 20.965 ;
        RECT 31.305 15.355 31.475 15.525 ;
        RECT 31.305 9.915 31.475 10.085 ;
        RECT 31.765 58.875 31.935 59.045 ;
        RECT 31.765 53.435 31.935 53.605 ;
        RECT 31.765 47.995 31.935 48.165 ;
        RECT 31.765 42.555 31.935 42.725 ;
        RECT 31.765 37.115 31.935 37.285 ;
        RECT 31.765 31.675 31.935 31.845 ;
        RECT 31.765 26.235 31.935 26.405 ;
        RECT 31.765 20.795 31.935 20.965 ;
        RECT 31.765 15.355 31.935 15.525 ;
        RECT 31.765 9.915 31.935 10.085 ;
        RECT 32.225 58.875 32.395 59.045 ;
        RECT 32.225 53.435 32.395 53.605 ;
        RECT 32.225 47.995 32.395 48.165 ;
        RECT 32.225 42.555 32.395 42.725 ;
        RECT 32.225 37.115 32.395 37.285 ;
        RECT 32.225 31.675 32.395 31.845 ;
        RECT 32.225 26.235 32.395 26.405 ;
        RECT 32.225 20.795 32.395 20.965 ;
        RECT 32.225 15.355 32.395 15.525 ;
        RECT 32.225 9.915 32.395 10.085 ;
        RECT 32.685 58.875 32.855 59.045 ;
        RECT 32.685 53.435 32.855 53.605 ;
        RECT 32.685 47.995 32.855 48.165 ;
        RECT 32.685 42.555 32.855 42.725 ;
        RECT 32.685 37.115 32.855 37.285 ;
        RECT 32.685 31.675 32.855 31.845 ;
        RECT 32.685 26.235 32.855 26.405 ;
        RECT 32.685 20.795 32.855 20.965 ;
        RECT 32.685 15.355 32.855 15.525 ;
        RECT 32.685 9.915 32.855 10.085 ;
        RECT 33.145 58.875 33.315 59.045 ;
        RECT 33.145 53.435 33.315 53.605 ;
        RECT 33.145 47.995 33.315 48.165 ;
        RECT 33.145 42.555 33.315 42.725 ;
        RECT 33.145 37.115 33.315 37.285 ;
        RECT 33.145 31.675 33.315 31.845 ;
        RECT 33.145 26.235 33.315 26.405 ;
        RECT 33.145 20.795 33.315 20.965 ;
        RECT 33.145 15.355 33.315 15.525 ;
        RECT 33.145 9.915 33.315 10.085 ;
        RECT 33.605 58.875 33.775 59.045 ;
        RECT 33.605 53.435 33.775 53.605 ;
        RECT 33.605 47.995 33.775 48.165 ;
        RECT 33.605 42.555 33.775 42.725 ;
        RECT 33.605 37.115 33.775 37.285 ;
        RECT 33.605 31.675 33.775 31.845 ;
        RECT 33.605 26.235 33.775 26.405 ;
        RECT 33.605 20.795 33.775 20.965 ;
        RECT 33.605 15.355 33.775 15.525 ;
        RECT 33.605 9.915 33.775 10.085 ;
        RECT 34.065 58.875 34.235 59.045 ;
        RECT 34.065 53.435 34.235 53.605 ;
        RECT 34.065 47.995 34.235 48.165 ;
        RECT 34.065 42.555 34.235 42.725 ;
        RECT 34.065 37.115 34.235 37.285 ;
        RECT 34.065 31.675 34.235 31.845 ;
        RECT 34.065 26.235 34.235 26.405 ;
        RECT 34.065 20.795 34.235 20.965 ;
        RECT 34.065 15.355 34.235 15.525 ;
        RECT 34.065 9.915 34.235 10.085 ;
        RECT 34.525 58.875 34.695 59.045 ;
        RECT 34.525 53.435 34.695 53.605 ;
        RECT 34.525 47.995 34.695 48.165 ;
        RECT 34.525 42.555 34.695 42.725 ;
        RECT 34.525 37.115 34.695 37.285 ;
        RECT 34.525 31.675 34.695 31.845 ;
        RECT 34.525 26.235 34.695 26.405 ;
        RECT 34.525 20.795 34.695 20.965 ;
        RECT 34.525 15.355 34.695 15.525 ;
        RECT 34.525 9.915 34.695 10.085 ;
        RECT 34.985 58.875 35.155 59.045 ;
        RECT 34.985 53.435 35.155 53.605 ;
        RECT 34.985 47.995 35.155 48.165 ;
        RECT 34.985 42.555 35.155 42.725 ;
        RECT 34.985 37.115 35.155 37.285 ;
        RECT 34.985 31.675 35.155 31.845 ;
        RECT 34.985 26.235 35.155 26.405 ;
        RECT 34.985 20.795 35.155 20.965 ;
        RECT 34.985 15.355 35.155 15.525 ;
        RECT 34.985 9.915 35.155 10.085 ;
        RECT 35.445 58.875 35.615 59.045 ;
        RECT 35.445 53.435 35.615 53.605 ;
        RECT 35.445 47.995 35.615 48.165 ;
        RECT 35.445 42.555 35.615 42.725 ;
        RECT 35.445 37.115 35.615 37.285 ;
        RECT 35.445 31.675 35.615 31.845 ;
        RECT 35.445 26.235 35.615 26.405 ;
        RECT 35.445 20.795 35.615 20.965 ;
        RECT 35.445 15.355 35.615 15.525 ;
        RECT 35.445 9.915 35.615 10.085 ;
        RECT 35.905 58.875 36.075 59.045 ;
        RECT 35.905 53.435 36.075 53.605 ;
        RECT 35.905 47.995 36.075 48.165 ;
        RECT 35.905 42.555 36.075 42.725 ;
        RECT 35.905 37.115 36.075 37.285 ;
        RECT 35.905 31.675 36.075 31.845 ;
        RECT 35.905 26.235 36.075 26.405 ;
        RECT 35.905 20.795 36.075 20.965 ;
        RECT 35.905 15.355 36.075 15.525 ;
        RECT 35.905 9.915 36.075 10.085 ;
        RECT 36.365 58.875 36.535 59.045 ;
        RECT 36.365 53.435 36.535 53.605 ;
        RECT 36.365 47.995 36.535 48.165 ;
        RECT 36.365 42.555 36.535 42.725 ;
        RECT 36.365 37.115 36.535 37.285 ;
        RECT 36.365 31.675 36.535 31.845 ;
        RECT 36.365 26.235 36.535 26.405 ;
        RECT 36.365 20.795 36.535 20.965 ;
        RECT 36.365 15.355 36.535 15.525 ;
        RECT 36.365 9.915 36.535 10.085 ;
        RECT 36.825 58.875 36.995 59.045 ;
        RECT 36.825 53.435 36.995 53.605 ;
        RECT 36.825 47.995 36.995 48.165 ;
        RECT 36.825 42.555 36.995 42.725 ;
        RECT 36.825 37.115 36.995 37.285 ;
        RECT 36.825 31.675 36.995 31.845 ;
        RECT 36.825 26.235 36.995 26.405 ;
        RECT 36.825 20.795 36.995 20.965 ;
        RECT 36.825 15.355 36.995 15.525 ;
        RECT 36.825 9.915 36.995 10.085 ;
        RECT 37.285 58.875 37.455 59.045 ;
        RECT 37.285 53.435 37.455 53.605 ;
        RECT 37.285 47.995 37.455 48.165 ;
        RECT 37.285 42.555 37.455 42.725 ;
        RECT 37.285 37.115 37.455 37.285 ;
        RECT 37.285 31.675 37.455 31.845 ;
        RECT 37.285 26.235 37.455 26.405 ;
        RECT 37.285 20.795 37.455 20.965 ;
        RECT 37.285 15.355 37.455 15.525 ;
        RECT 37.285 9.915 37.455 10.085 ;
        RECT 37.745 58.875 37.915 59.045 ;
        RECT 37.745 53.435 37.915 53.605 ;
        RECT 37.745 47.995 37.915 48.165 ;
        RECT 37.745 42.555 37.915 42.725 ;
        RECT 37.745 37.115 37.915 37.285 ;
        RECT 37.745 31.675 37.915 31.845 ;
        RECT 37.745 26.235 37.915 26.405 ;
        RECT 37.745 20.795 37.915 20.965 ;
        RECT 37.745 15.355 37.915 15.525 ;
        RECT 37.745 9.915 37.915 10.085 ;
        RECT 38.205 58.875 38.375 59.045 ;
        RECT 38.205 53.435 38.375 53.605 ;
        RECT 38.205 47.995 38.375 48.165 ;
        RECT 38.205 42.555 38.375 42.725 ;
        RECT 38.205 37.115 38.375 37.285 ;
        RECT 38.205 31.675 38.375 31.845 ;
        RECT 38.205 26.235 38.375 26.405 ;
        RECT 38.205 20.795 38.375 20.965 ;
        RECT 38.205 15.355 38.375 15.525 ;
        RECT 38.205 9.915 38.375 10.085 ;
        RECT 38.665 58.875 38.835 59.045 ;
        RECT 38.665 53.435 38.835 53.605 ;
        RECT 38.665 47.995 38.835 48.165 ;
        RECT 38.665 42.555 38.835 42.725 ;
        RECT 38.665 37.115 38.835 37.285 ;
        RECT 38.665 31.675 38.835 31.845 ;
        RECT 38.665 26.235 38.835 26.405 ;
        RECT 38.665 20.795 38.835 20.965 ;
        RECT 38.665 15.355 38.835 15.525 ;
        RECT 38.665 9.915 38.835 10.085 ;
        RECT 39.125 58.875 39.295 59.045 ;
        RECT 39.125 53.435 39.295 53.605 ;
        RECT 39.125 47.995 39.295 48.165 ;
        RECT 39.125 42.555 39.295 42.725 ;
        RECT 39.125 37.115 39.295 37.285 ;
        RECT 39.125 31.675 39.295 31.845 ;
        RECT 39.125 26.235 39.295 26.405 ;
        RECT 39.125 20.795 39.295 20.965 ;
        RECT 39.125 15.355 39.295 15.525 ;
        RECT 39.125 9.915 39.295 10.085 ;
        RECT 39.585 58.875 39.755 59.045 ;
        RECT 39.585 53.435 39.755 53.605 ;
        RECT 39.585 47.995 39.755 48.165 ;
        RECT 39.585 42.555 39.755 42.725 ;
        RECT 39.585 37.115 39.755 37.285 ;
        RECT 39.585 31.675 39.755 31.845 ;
        RECT 39.585 26.235 39.755 26.405 ;
        RECT 39.585 20.795 39.755 20.965 ;
        RECT 39.585 15.355 39.755 15.525 ;
        RECT 39.585 9.915 39.755 10.085 ;
        RECT 40.045 58.875 40.215 59.045 ;
        RECT 40.045 53.435 40.215 53.605 ;
        RECT 40.045 47.995 40.215 48.165 ;
        RECT 40.045 42.555 40.215 42.725 ;
        RECT 40.045 37.115 40.215 37.285 ;
        RECT 40.045 31.675 40.215 31.845 ;
        RECT 40.045 26.235 40.215 26.405 ;
        RECT 40.045 20.795 40.215 20.965 ;
        RECT 40.045 15.355 40.215 15.525 ;
        RECT 40.045 9.915 40.215 10.085 ;
        RECT 40.505 58.875 40.675 59.045 ;
        RECT 40.505 53.435 40.675 53.605 ;
        RECT 40.505 47.995 40.675 48.165 ;
        RECT 40.505 42.555 40.675 42.725 ;
        RECT 40.505 37.115 40.675 37.285 ;
        RECT 40.505 31.675 40.675 31.845 ;
        RECT 40.505 26.235 40.675 26.405 ;
        RECT 40.505 20.795 40.675 20.965 ;
        RECT 40.505 15.355 40.675 15.525 ;
        RECT 40.505 9.915 40.675 10.085 ;
        RECT 40.965 58.875 41.135 59.045 ;
        RECT 40.965 53.435 41.135 53.605 ;
        RECT 40.965 47.995 41.135 48.165 ;
        RECT 40.965 42.555 41.135 42.725 ;
        RECT 40.965 37.115 41.135 37.285 ;
        RECT 40.965 31.675 41.135 31.845 ;
        RECT 40.965 26.235 41.135 26.405 ;
        RECT 40.965 20.795 41.135 20.965 ;
        RECT 40.965 15.355 41.135 15.525 ;
        RECT 40.965 9.915 41.135 10.085 ;
        RECT 41.425 58.875 41.595 59.045 ;
        RECT 41.425 53.435 41.595 53.605 ;
        RECT 41.425 47.995 41.595 48.165 ;
        RECT 41.425 42.555 41.595 42.725 ;
        RECT 41.425 37.115 41.595 37.285 ;
        RECT 41.425 31.675 41.595 31.845 ;
        RECT 41.425 26.235 41.595 26.405 ;
        RECT 41.425 20.795 41.595 20.965 ;
        RECT 41.425 15.355 41.595 15.525 ;
        RECT 41.425 9.915 41.595 10.085 ;
        RECT 41.885 58.875 42.055 59.045 ;
        RECT 41.885 53.435 42.055 53.605 ;
        RECT 41.885 47.995 42.055 48.165 ;
        RECT 41.885 42.555 42.055 42.725 ;
        RECT 41.885 37.115 42.055 37.285 ;
        RECT 41.885 31.675 42.055 31.845 ;
        RECT 41.885 26.235 42.055 26.405 ;
        RECT 41.885 20.795 42.055 20.965 ;
        RECT 41.885 15.355 42.055 15.525 ;
        RECT 41.885 9.915 42.055 10.085 ;
        RECT 42.345 58.875 42.515 59.045 ;
        RECT 42.345 53.435 42.515 53.605 ;
        RECT 42.345 47.995 42.515 48.165 ;
        RECT 42.345 42.555 42.515 42.725 ;
        RECT 42.345 37.115 42.515 37.285 ;
        RECT 42.345 31.675 42.515 31.845 ;
        RECT 42.345 26.235 42.515 26.405 ;
        RECT 42.345 20.795 42.515 20.965 ;
        RECT 42.345 15.355 42.515 15.525 ;
        RECT 42.345 9.915 42.515 10.085 ;
        RECT 42.805 58.875 42.975 59.045 ;
        RECT 42.805 53.435 42.975 53.605 ;
        RECT 42.805 47.995 42.975 48.165 ;
        RECT 42.805 42.555 42.975 42.725 ;
        RECT 42.805 37.115 42.975 37.285 ;
        RECT 42.805 31.675 42.975 31.845 ;
        RECT 42.805 26.235 42.975 26.405 ;
        RECT 42.805 20.795 42.975 20.965 ;
        RECT 42.805 15.355 42.975 15.525 ;
        RECT 42.805 9.915 42.975 10.085 ;
        RECT 43.265 58.875 43.435 59.045 ;
        RECT 43.265 53.435 43.435 53.605 ;
        RECT 43.265 47.995 43.435 48.165 ;
        RECT 43.265 42.555 43.435 42.725 ;
        RECT 43.265 37.115 43.435 37.285 ;
        RECT 43.265 31.675 43.435 31.845 ;
        RECT 43.265 26.235 43.435 26.405 ;
        RECT 43.265 20.795 43.435 20.965 ;
        RECT 43.265 15.355 43.435 15.525 ;
        RECT 43.265 9.915 43.435 10.085 ;
        RECT 43.725 58.875 43.895 59.045 ;
        RECT 43.725 53.435 43.895 53.605 ;
        RECT 43.725 47.995 43.895 48.165 ;
        RECT 43.725 42.555 43.895 42.725 ;
        RECT 43.725 37.115 43.895 37.285 ;
        RECT 43.725 31.675 43.895 31.845 ;
        RECT 43.725 26.235 43.895 26.405 ;
        RECT 43.725 20.795 43.895 20.965 ;
        RECT 43.725 15.355 43.895 15.525 ;
        RECT 43.725 9.915 43.895 10.085 ;
        RECT 44.185 58.875 44.355 59.045 ;
        RECT 44.185 53.435 44.355 53.605 ;
        RECT 44.185 47.995 44.355 48.165 ;
        RECT 44.185 42.555 44.355 42.725 ;
        RECT 44.185 37.115 44.355 37.285 ;
        RECT 44.185 31.675 44.355 31.845 ;
        RECT 44.185 26.235 44.355 26.405 ;
        RECT 44.185 20.795 44.355 20.965 ;
        RECT 44.185 15.355 44.355 15.525 ;
        RECT 44.185 9.915 44.355 10.085 ;
        RECT 44.645 58.875 44.815 59.045 ;
        RECT 44.645 53.435 44.815 53.605 ;
        RECT 44.645 47.995 44.815 48.165 ;
        RECT 44.645 42.555 44.815 42.725 ;
        RECT 44.645 37.115 44.815 37.285 ;
        RECT 44.645 31.675 44.815 31.845 ;
        RECT 44.645 26.235 44.815 26.405 ;
        RECT 44.645 20.795 44.815 20.965 ;
        RECT 44.645 15.355 44.815 15.525 ;
        RECT 44.645 9.915 44.815 10.085 ;
        RECT 45.105 58.875 45.275 59.045 ;
        RECT 45.105 53.435 45.275 53.605 ;
        RECT 45.105 47.995 45.275 48.165 ;
        RECT 45.105 42.555 45.275 42.725 ;
        RECT 45.105 37.115 45.275 37.285 ;
        RECT 45.105 31.675 45.275 31.845 ;
        RECT 45.105 26.235 45.275 26.405 ;
        RECT 45.105 20.795 45.275 20.965 ;
        RECT 45.105 15.355 45.275 15.525 ;
        RECT 45.105 9.915 45.275 10.085 ;
        RECT 45.565 58.875 45.735 59.045 ;
        RECT 45.565 53.435 45.735 53.605 ;
        RECT 45.565 47.995 45.735 48.165 ;
        RECT 45.565 42.555 45.735 42.725 ;
        RECT 45.565 37.115 45.735 37.285 ;
        RECT 45.565 31.675 45.735 31.845 ;
        RECT 45.565 26.235 45.735 26.405 ;
        RECT 45.565 20.795 45.735 20.965 ;
        RECT 45.565 15.355 45.735 15.525 ;
        RECT 45.565 9.915 45.735 10.085 ;
        RECT 46.025 58.875 46.195 59.045 ;
        RECT 46.025 53.435 46.195 53.605 ;
        RECT 46.025 47.995 46.195 48.165 ;
        RECT 46.025 42.555 46.195 42.725 ;
        RECT 46.025 37.115 46.195 37.285 ;
        RECT 46.025 31.675 46.195 31.845 ;
        RECT 46.025 26.235 46.195 26.405 ;
        RECT 46.025 20.795 46.195 20.965 ;
        RECT 46.025 15.355 46.195 15.525 ;
        RECT 46.025 9.915 46.195 10.085 ;
        RECT 46.485 58.875 46.655 59.045 ;
        RECT 46.485 53.435 46.655 53.605 ;
        RECT 46.485 47.995 46.655 48.165 ;
        RECT 46.485 42.555 46.655 42.725 ;
        RECT 46.485 37.115 46.655 37.285 ;
        RECT 46.485 31.675 46.655 31.845 ;
        RECT 46.485 26.235 46.655 26.405 ;
        RECT 46.485 20.795 46.655 20.965 ;
        RECT 46.485 15.355 46.655 15.525 ;
        RECT 46.485 9.915 46.655 10.085 ;
        RECT 46.945 58.875 47.115 59.045 ;
        RECT 46.945 53.435 47.115 53.605 ;
        RECT 46.945 47.995 47.115 48.165 ;
        RECT 46.945 42.555 47.115 42.725 ;
        RECT 46.945 37.115 47.115 37.285 ;
        RECT 46.945 31.675 47.115 31.845 ;
        RECT 46.945 26.235 47.115 26.405 ;
        RECT 46.945 20.795 47.115 20.965 ;
        RECT 46.945 15.355 47.115 15.525 ;
        RECT 46.945 9.915 47.115 10.085 ;
        RECT 47.405 58.875 47.575 59.045 ;
        RECT 47.405 53.435 47.575 53.605 ;
        RECT 47.405 47.995 47.575 48.165 ;
        RECT 47.405 42.555 47.575 42.725 ;
        RECT 47.405 37.115 47.575 37.285 ;
        RECT 47.405 31.675 47.575 31.845 ;
        RECT 47.405 26.235 47.575 26.405 ;
        RECT 47.405 20.795 47.575 20.965 ;
        RECT 47.405 15.355 47.575 15.525 ;
        RECT 47.405 9.915 47.575 10.085 ;
        RECT 47.865 58.875 48.035 59.045 ;
        RECT 47.865 53.435 48.035 53.605 ;
        RECT 47.865 47.995 48.035 48.165 ;
        RECT 47.865 42.555 48.035 42.725 ;
        RECT 47.865 37.115 48.035 37.285 ;
        RECT 47.865 31.675 48.035 31.845 ;
        RECT 47.865 26.235 48.035 26.405 ;
        RECT 47.865 20.795 48.035 20.965 ;
        RECT 47.865 15.355 48.035 15.525 ;
        RECT 47.865 9.915 48.035 10.085 ;
        RECT 48.325 58.875 48.495 59.045 ;
        RECT 48.325 53.435 48.495 53.605 ;
        RECT 48.325 47.995 48.495 48.165 ;
        RECT 48.325 42.555 48.495 42.725 ;
        RECT 48.325 37.115 48.495 37.285 ;
        RECT 48.325 31.675 48.495 31.845 ;
        RECT 48.325 26.235 48.495 26.405 ;
        RECT 48.325 20.795 48.495 20.965 ;
        RECT 48.325 15.355 48.495 15.525 ;
        RECT 48.325 9.915 48.495 10.085 ;
        RECT 48.785 58.875 48.955 59.045 ;
        RECT 48.785 53.435 48.955 53.605 ;
        RECT 48.785 47.995 48.955 48.165 ;
        RECT 48.785 42.555 48.955 42.725 ;
        RECT 48.785 37.115 48.955 37.285 ;
        RECT 48.785 31.675 48.955 31.845 ;
        RECT 48.785 26.235 48.955 26.405 ;
        RECT 48.785 20.795 48.955 20.965 ;
        RECT 48.785 15.355 48.955 15.525 ;
        RECT 48.785 9.915 48.955 10.085 ;
        RECT 49.245 58.875 49.415 59.045 ;
        RECT 49.245 53.435 49.415 53.605 ;
        RECT 49.245 47.995 49.415 48.165 ;
        RECT 49.245 42.555 49.415 42.725 ;
        RECT 49.245 37.115 49.415 37.285 ;
        RECT 49.245 31.675 49.415 31.845 ;
        RECT 49.245 26.235 49.415 26.405 ;
        RECT 49.245 20.795 49.415 20.965 ;
        RECT 49.245 15.355 49.415 15.525 ;
        RECT 49.245 9.915 49.415 10.085 ;
        RECT 49.705 58.875 49.875 59.045 ;
        RECT 49.705 53.435 49.875 53.605 ;
        RECT 49.705 47.995 49.875 48.165 ;
        RECT 49.705 42.555 49.875 42.725 ;
        RECT 49.705 37.115 49.875 37.285 ;
        RECT 49.705 31.675 49.875 31.845 ;
        RECT 49.705 26.235 49.875 26.405 ;
        RECT 49.705 20.795 49.875 20.965 ;
        RECT 49.705 15.355 49.875 15.525 ;
        RECT 49.705 9.915 49.875 10.085 ;
        RECT 50.165 58.875 50.335 59.045 ;
        RECT 50.165 53.435 50.335 53.605 ;
        RECT 50.165 47.995 50.335 48.165 ;
        RECT 50.165 42.555 50.335 42.725 ;
        RECT 50.165 37.115 50.335 37.285 ;
        RECT 50.165 31.675 50.335 31.845 ;
        RECT 50.165 26.235 50.335 26.405 ;
        RECT 50.165 20.795 50.335 20.965 ;
        RECT 50.165 15.355 50.335 15.525 ;
        RECT 50.165 9.915 50.335 10.085 ;
        RECT 50.625 58.875 50.795 59.045 ;
        RECT 50.625 53.435 50.795 53.605 ;
        RECT 50.625 47.995 50.795 48.165 ;
        RECT 50.625 42.555 50.795 42.725 ;
        RECT 50.625 37.115 50.795 37.285 ;
        RECT 50.625 31.675 50.795 31.845 ;
        RECT 50.625 26.235 50.795 26.405 ;
        RECT 50.625 20.795 50.795 20.965 ;
        RECT 50.625 15.355 50.795 15.525 ;
        RECT 50.625 9.915 50.795 10.085 ;
        RECT 51.085 58.875 51.255 59.045 ;
        RECT 51.085 53.435 51.255 53.605 ;
        RECT 51.085 47.995 51.255 48.165 ;
        RECT 51.085 42.555 51.255 42.725 ;
        RECT 51.085 37.115 51.255 37.285 ;
        RECT 51.085 31.675 51.255 31.845 ;
        RECT 51.085 26.235 51.255 26.405 ;
        RECT 51.085 20.795 51.255 20.965 ;
        RECT 51.085 15.355 51.255 15.525 ;
        RECT 51.085 9.915 51.255 10.085 ;
        RECT 51.545 58.875 51.715 59.045 ;
        RECT 51.545 53.435 51.715 53.605 ;
        RECT 51.545 47.995 51.715 48.165 ;
        RECT 51.545 42.555 51.715 42.725 ;
        RECT 51.545 37.115 51.715 37.285 ;
        RECT 51.545 31.675 51.715 31.845 ;
        RECT 51.545 26.235 51.715 26.405 ;
        RECT 51.545 20.795 51.715 20.965 ;
        RECT 51.545 15.355 51.715 15.525 ;
        RECT 51.545 9.915 51.715 10.085 ;
        RECT 52.005 58.875 52.175 59.045 ;
        RECT 52.005 53.435 52.175 53.605 ;
        RECT 52.005 47.995 52.175 48.165 ;
        RECT 52.005 42.555 52.175 42.725 ;
        RECT 52.005 37.115 52.175 37.285 ;
        RECT 52.005 31.675 52.175 31.845 ;
        RECT 52.005 26.235 52.175 26.405 ;
        RECT 52.005 20.795 52.175 20.965 ;
        RECT 52.005 15.355 52.175 15.525 ;
        RECT 52.005 9.915 52.175 10.085 ;
        RECT 52.465 58.875 52.635 59.045 ;
        RECT 52.465 53.435 52.635 53.605 ;
        RECT 52.465 47.995 52.635 48.165 ;
        RECT 52.465 42.555 52.635 42.725 ;
        RECT 52.465 37.115 52.635 37.285 ;
        RECT 52.465 31.675 52.635 31.845 ;
        RECT 52.465 26.235 52.635 26.405 ;
        RECT 52.465 20.795 52.635 20.965 ;
        RECT 52.465 15.355 52.635 15.525 ;
        RECT 52.465 9.915 52.635 10.085 ;
        RECT 52.925 58.875 53.095 59.045 ;
        RECT 52.925 53.435 53.095 53.605 ;
        RECT 52.925 47.995 53.095 48.165 ;
        RECT 52.925 42.555 53.095 42.725 ;
        RECT 52.925 37.115 53.095 37.285 ;
        RECT 52.925 31.675 53.095 31.845 ;
        RECT 52.925 26.235 53.095 26.405 ;
        RECT 52.925 20.795 53.095 20.965 ;
        RECT 52.925 15.355 53.095 15.525 ;
        RECT 52.925 9.915 53.095 10.085 ;
        RECT 53.385 58.875 53.555 59.045 ;
        RECT 53.385 53.435 53.555 53.605 ;
        RECT 53.385 47.995 53.555 48.165 ;
        RECT 53.385 42.555 53.555 42.725 ;
        RECT 53.385 37.115 53.555 37.285 ;
        RECT 53.385 31.675 53.555 31.845 ;
        RECT 53.385 26.235 53.555 26.405 ;
        RECT 53.385 20.795 53.555 20.965 ;
        RECT 53.385 15.355 53.555 15.525 ;
        RECT 53.385 9.915 53.555 10.085 ;
        RECT 53.845 58.875 54.015 59.045 ;
        RECT 53.845 53.435 54.015 53.605 ;
        RECT 53.845 47.995 54.015 48.165 ;
        RECT 53.845 42.555 54.015 42.725 ;
        RECT 53.845 37.115 54.015 37.285 ;
        RECT 53.845 31.675 54.015 31.845 ;
        RECT 53.845 26.235 54.015 26.405 ;
        RECT 53.845 20.795 54.015 20.965 ;
        RECT 53.845 15.355 54.015 15.525 ;
        RECT 53.845 9.915 54.015 10.085 ;
        RECT 54.305 58.875 54.475 59.045 ;
        RECT 54.305 53.435 54.475 53.605 ;
        RECT 54.305 47.995 54.475 48.165 ;
        RECT 54.305 42.555 54.475 42.725 ;
        RECT 54.305 37.115 54.475 37.285 ;
        RECT 54.305 31.675 54.475 31.845 ;
        RECT 54.305 26.235 54.475 26.405 ;
        RECT 54.305 20.795 54.475 20.965 ;
        RECT 54.305 15.355 54.475 15.525 ;
        RECT 54.305 9.915 54.475 10.085 ;
        RECT 54.765 58.875 54.935 59.045 ;
        RECT 54.765 53.435 54.935 53.605 ;
        RECT 54.765 47.995 54.935 48.165 ;
        RECT 54.765 42.555 54.935 42.725 ;
        RECT 54.765 37.115 54.935 37.285 ;
        RECT 54.765 31.675 54.935 31.845 ;
        RECT 54.765 26.235 54.935 26.405 ;
        RECT 54.765 20.795 54.935 20.965 ;
        RECT 54.765 15.355 54.935 15.525 ;
        RECT 54.765 9.915 54.935 10.085 ;
        RECT 55.225 58.875 55.395 59.045 ;
        RECT 55.225 53.435 55.395 53.605 ;
        RECT 55.225 47.995 55.395 48.165 ;
        RECT 55.225 42.555 55.395 42.725 ;
        RECT 55.225 37.115 55.395 37.285 ;
        RECT 55.225 31.675 55.395 31.845 ;
        RECT 55.225 26.235 55.395 26.405 ;
        RECT 55.225 20.795 55.395 20.965 ;
        RECT 55.225 15.355 55.395 15.525 ;
        RECT 55.225 9.915 55.395 10.085 ;
        RECT 55.685 58.875 55.855 59.045 ;
        RECT 55.685 53.435 55.855 53.605 ;
        RECT 55.685 47.995 55.855 48.165 ;
        RECT 55.685 42.555 55.855 42.725 ;
        RECT 55.685 37.115 55.855 37.285 ;
        RECT 55.685 31.675 55.855 31.845 ;
        RECT 55.685 26.235 55.855 26.405 ;
        RECT 55.685 20.795 55.855 20.965 ;
        RECT 55.685 15.355 55.855 15.525 ;
        RECT 55.685 9.915 55.855 10.085 ;
      LAYER via2 ;
        RECT 11.97 57.84 12.17 58.04 ;
        RECT 11.97 53.76 12.17 53.96 ;
        RECT 11.97 49.68 12.17 49.88 ;
        RECT 11.97 45.6 12.17 45.8 ;
        RECT 11.97 41.52 12.17 41.72 ;
        RECT 11.97 37.44 12.17 37.64 ;
        RECT 11.97 33.36 12.17 33.56 ;
        RECT 11.97 29.28 12.17 29.48 ;
        RECT 11.97 25.2 12.17 25.4 ;
        RECT 11.97 21.12 12.17 21.32 ;
        RECT 11.97 17.04 12.17 17.24 ;
        RECT 11.97 12.96 12.17 13.16 ;
        RECT 14.73 57.84 14.93 58.04 ;
        RECT 14.73 53.76 14.93 53.96 ;
        RECT 14.73 49.68 14.93 49.88 ;
        RECT 14.73 45.6 14.93 45.8 ;
        RECT 14.73 41.52 14.93 41.72 ;
        RECT 14.73 37.44 14.93 37.64 ;
        RECT 14.73 33.36 14.93 33.56 ;
        RECT 14.73 29.28 14.93 29.48 ;
        RECT 14.73 25.2 14.93 25.4 ;
        RECT 14.73 21.12 14.93 21.32 ;
        RECT 14.73 17.04 14.93 17.24 ;
        RECT 14.73 12.96 14.93 13.16 ;
        RECT 17.49 57.84 17.69 58.04 ;
        RECT 17.49 53.76 17.69 53.96 ;
        RECT 17.49 49.68 17.69 49.88 ;
        RECT 17.49 45.6 17.69 45.8 ;
        RECT 17.49 41.52 17.69 41.72 ;
        RECT 17.49 37.44 17.69 37.64 ;
        RECT 17.49 33.36 17.69 33.56 ;
        RECT 17.49 29.28 17.69 29.48 ;
        RECT 17.49 25.2 17.69 25.4 ;
        RECT 17.49 21.12 17.69 21.32 ;
        RECT 17.49 17.04 17.69 17.24 ;
        RECT 17.49 12.96 17.69 13.16 ;
        RECT 20.25 57.84 20.45 58.04 ;
        RECT 20.25 53.76 20.45 53.96 ;
        RECT 20.25 49.68 20.45 49.88 ;
        RECT 20.25 45.6 20.45 45.8 ;
        RECT 20.25 41.52 20.45 41.72 ;
        RECT 20.25 37.44 20.45 37.64 ;
        RECT 20.25 33.36 20.45 33.56 ;
        RECT 20.25 29.28 20.45 29.48 ;
        RECT 20.25 25.2 20.45 25.4 ;
        RECT 20.25 21.12 20.45 21.32 ;
        RECT 20.25 17.04 20.45 17.24 ;
        RECT 20.25 12.96 20.45 13.16 ;
        RECT 23.01 57.84 23.21 58.04 ;
        RECT 23.01 53.76 23.21 53.96 ;
        RECT 23.01 49.68 23.21 49.88 ;
        RECT 23.01 45.6 23.21 45.8 ;
        RECT 23.01 41.52 23.21 41.72 ;
        RECT 23.01 37.44 23.21 37.64 ;
        RECT 23.01 33.36 23.21 33.56 ;
        RECT 23.01 29.28 23.21 29.48 ;
        RECT 23.01 25.2 23.21 25.4 ;
        RECT 23.01 21.12 23.21 21.32 ;
        RECT 23.01 17.04 23.21 17.24 ;
        RECT 23.01 12.96 23.21 13.16 ;
        RECT 25.77 57.84 25.97 58.04 ;
        RECT 25.77 53.76 25.97 53.96 ;
        RECT 25.77 49.68 25.97 49.88 ;
        RECT 25.77 45.6 25.97 45.8 ;
        RECT 25.77 41.52 25.97 41.72 ;
        RECT 25.77 37.44 25.97 37.64 ;
        RECT 25.77 33.36 25.97 33.56 ;
        RECT 25.77 29.28 25.97 29.48 ;
        RECT 25.77 25.2 25.97 25.4 ;
        RECT 25.77 21.12 25.97 21.32 ;
        RECT 25.77 17.04 25.97 17.24 ;
        RECT 25.77 12.96 25.97 13.16 ;
        RECT 28.53 57.84 28.73 58.04 ;
        RECT 28.53 53.76 28.73 53.96 ;
        RECT 28.53 49.68 28.73 49.88 ;
        RECT 28.53 45.6 28.73 45.8 ;
        RECT 28.53 41.52 28.73 41.72 ;
        RECT 28.53 37.44 28.73 37.64 ;
        RECT 28.53 33.36 28.73 33.56 ;
        RECT 28.53 29.28 28.73 29.48 ;
        RECT 28.53 25.2 28.73 25.4 ;
        RECT 28.53 21.12 28.73 21.32 ;
        RECT 28.53 17.04 28.73 17.24 ;
        RECT 28.53 12.96 28.73 13.16 ;
        RECT 31.29 57.84 31.49 58.04 ;
        RECT 31.29 53.76 31.49 53.96 ;
        RECT 31.29 49.68 31.49 49.88 ;
        RECT 31.29 45.6 31.49 45.8 ;
        RECT 31.29 41.52 31.49 41.72 ;
        RECT 31.29 37.44 31.49 37.64 ;
        RECT 31.29 33.36 31.49 33.56 ;
        RECT 31.29 29.28 31.49 29.48 ;
        RECT 31.29 25.2 31.49 25.4 ;
        RECT 31.29 21.12 31.49 21.32 ;
        RECT 31.29 17.04 31.49 17.24 ;
        RECT 31.29 12.96 31.49 13.16 ;
        RECT 34.05 57.84 34.25 58.04 ;
        RECT 34.05 53.76 34.25 53.96 ;
        RECT 34.05 49.68 34.25 49.88 ;
        RECT 34.05 45.6 34.25 45.8 ;
        RECT 34.05 41.52 34.25 41.72 ;
        RECT 34.05 37.44 34.25 37.64 ;
        RECT 34.05 33.36 34.25 33.56 ;
        RECT 34.05 29.28 34.25 29.48 ;
        RECT 34.05 25.2 34.25 25.4 ;
        RECT 34.05 21.12 34.25 21.32 ;
        RECT 34.05 17.04 34.25 17.24 ;
        RECT 34.05 12.96 34.25 13.16 ;
        RECT 36.81 57.84 37.01 58.04 ;
        RECT 36.81 53.76 37.01 53.96 ;
        RECT 36.81 49.68 37.01 49.88 ;
        RECT 36.81 45.6 37.01 45.8 ;
        RECT 36.81 41.52 37.01 41.72 ;
        RECT 36.81 37.44 37.01 37.64 ;
        RECT 36.81 33.36 37.01 33.56 ;
        RECT 36.81 29.28 37.01 29.48 ;
        RECT 36.81 25.2 37.01 25.4 ;
        RECT 36.81 21.12 37.01 21.32 ;
        RECT 36.81 17.04 37.01 17.24 ;
        RECT 36.81 12.96 37.01 13.16 ;
        RECT 39.57 57.84 39.77 58.04 ;
        RECT 39.57 53.76 39.77 53.96 ;
        RECT 39.57 49.68 39.77 49.88 ;
        RECT 39.57 45.6 39.77 45.8 ;
        RECT 39.57 41.52 39.77 41.72 ;
        RECT 39.57 37.44 39.77 37.64 ;
        RECT 39.57 33.36 39.77 33.56 ;
        RECT 39.57 29.28 39.77 29.48 ;
        RECT 39.57 25.2 39.77 25.4 ;
        RECT 39.57 21.12 39.77 21.32 ;
        RECT 39.57 17.04 39.77 17.24 ;
        RECT 39.57 12.96 39.77 13.16 ;
        RECT 42.33 57.84 42.53 58.04 ;
        RECT 42.33 53.76 42.53 53.96 ;
        RECT 42.33 49.68 42.53 49.88 ;
        RECT 42.33 45.6 42.53 45.8 ;
        RECT 42.33 41.52 42.53 41.72 ;
        RECT 42.33 37.44 42.53 37.64 ;
        RECT 42.33 33.36 42.53 33.56 ;
        RECT 42.33 29.28 42.53 29.48 ;
        RECT 42.33 25.2 42.53 25.4 ;
        RECT 42.33 21.12 42.53 21.32 ;
        RECT 42.33 17.04 42.53 17.24 ;
        RECT 42.33 12.96 42.53 13.16 ;
        RECT 45.09 57.84 45.29 58.04 ;
        RECT 45.09 53.76 45.29 53.96 ;
        RECT 45.09 49.68 45.29 49.88 ;
        RECT 45.09 45.6 45.29 45.8 ;
        RECT 45.09 41.52 45.29 41.72 ;
        RECT 45.09 37.44 45.29 37.64 ;
        RECT 45.09 33.36 45.29 33.56 ;
        RECT 45.09 29.28 45.29 29.48 ;
        RECT 45.09 25.2 45.29 25.4 ;
        RECT 45.09 21.12 45.29 21.32 ;
        RECT 45.09 17.04 45.29 17.24 ;
        RECT 45.09 12.96 45.29 13.16 ;
        RECT 47.85 57.84 48.05 58.04 ;
        RECT 47.85 53.76 48.05 53.96 ;
        RECT 47.85 49.68 48.05 49.88 ;
        RECT 47.85 45.6 48.05 45.8 ;
        RECT 47.85 41.52 48.05 41.72 ;
        RECT 47.85 37.44 48.05 37.64 ;
        RECT 47.85 33.36 48.05 33.56 ;
        RECT 47.85 29.28 48.05 29.48 ;
        RECT 47.85 25.2 48.05 25.4 ;
        RECT 47.85 21.12 48.05 21.32 ;
        RECT 47.85 17.04 48.05 17.24 ;
        RECT 47.85 12.96 48.05 13.16 ;
        RECT 50.61 57.84 50.81 58.04 ;
        RECT 50.61 53.76 50.81 53.96 ;
        RECT 50.61 49.68 50.81 49.88 ;
        RECT 50.61 45.6 50.81 45.8 ;
        RECT 50.61 41.52 50.81 41.72 ;
        RECT 50.61 37.44 50.81 37.64 ;
        RECT 50.61 33.36 50.81 33.56 ;
        RECT 50.61 29.28 50.81 29.48 ;
        RECT 50.61 25.2 50.81 25.4 ;
        RECT 50.61 21.12 50.81 21.32 ;
        RECT 50.61 17.04 50.81 17.24 ;
        RECT 50.61 12.96 50.81 13.16 ;
        RECT 53.37 57.84 53.57 58.04 ;
        RECT 53.37 53.76 53.57 53.96 ;
        RECT 53.37 49.68 53.57 49.88 ;
        RECT 53.37 45.6 53.57 45.8 ;
        RECT 53.37 41.52 53.57 41.72 ;
        RECT 53.37 37.44 53.57 37.64 ;
        RECT 53.37 33.36 53.57 33.56 ;
        RECT 53.37 29.28 53.57 29.48 ;
        RECT 53.37 25.2 53.57 25.4 ;
        RECT 53.37 21.12 53.57 21.32 ;
        RECT 53.37 17.04 53.57 17.24 ;
        RECT 53.37 12.96 53.57 13.16 ;
        RECT 56.13 57.84 56.33 58.04 ;
        RECT 56.13 53.76 56.33 53.96 ;
        RECT 56.13 49.68 56.33 49.88 ;
        RECT 56.13 45.6 56.33 45.8 ;
        RECT 56.13 41.52 56.33 41.72 ;
        RECT 56.13 37.44 56.33 37.64 ;
        RECT 56.13 33.36 56.33 33.56 ;
        RECT 56.13 29.28 56.33 29.48 ;
        RECT 56.13 25.2 56.33 25.4 ;
        RECT 56.13 21.12 56.33 21.32 ;
        RECT 56.13 17.04 56.33 17.24 ;
        RECT 56.13 12.96 56.33 13.16 ;
        RECT 58.89 57.84 59.09 58.04 ;
        RECT 58.89 53.76 59.09 53.96 ;
        RECT 58.89 49.68 59.09 49.88 ;
        RECT 58.89 45.6 59.09 45.8 ;
        RECT 58.89 41.52 59.09 41.72 ;
        RECT 58.89 37.44 59.09 37.64 ;
        RECT 58.89 33.36 59.09 33.56 ;
        RECT 58.89 29.28 59.09 29.48 ;
        RECT 58.89 25.2 59.09 25.4 ;
        RECT 58.89 21.12 59.09 21.32 ;
        RECT 58.89 17.04 59.09 17.24 ;
        RECT 58.89 12.96 59.09 13.16 ;
        RECT 61.65 57.84 61.85 58.04 ;
        RECT 61.65 53.76 61.85 53.96 ;
        RECT 61.65 49.68 61.85 49.88 ;
        RECT 61.65 45.6 61.85 45.8 ;
        RECT 61.65 41.52 61.85 41.72 ;
        RECT 61.65 37.44 61.85 37.64 ;
        RECT 61.65 33.36 61.85 33.56 ;
        RECT 61.65 29.28 61.85 29.48 ;
        RECT 61.65 25.2 61.85 25.4 ;
        RECT 61.65 21.12 61.85 21.32 ;
        RECT 61.65 17.04 61.85 17.24 ;
        RECT 61.65 12.96 61.85 13.16 ;
        RECT 64.41 57.84 64.61 58.04 ;
        RECT 64.41 53.76 64.61 53.96 ;
        RECT 64.41 49.68 64.61 49.88 ;
        RECT 64.41 45.6 64.61 45.8 ;
        RECT 64.41 41.52 64.61 41.72 ;
        RECT 64.41 37.44 64.61 37.64 ;
        RECT 64.41 33.36 64.61 33.56 ;
        RECT 64.41 29.28 64.61 29.48 ;
        RECT 64.41 25.2 64.61 25.4 ;
        RECT 64.41 21.12 64.61 21.32 ;
        RECT 64.41 17.04 64.61 17.24 ;
        RECT 64.41 12.96 64.61 13.16 ;
        RECT 67.17 57.84 67.37 58.04 ;
        RECT 67.17 53.76 67.37 53.96 ;
        RECT 67.17 49.68 67.37 49.88 ;
        RECT 67.17 45.6 67.37 45.8 ;
        RECT 67.17 41.52 67.37 41.72 ;
        RECT 67.17 37.44 67.37 37.64 ;
        RECT 67.17 33.36 67.37 33.56 ;
        RECT 67.17 29.28 67.37 29.48 ;
        RECT 67.17 25.2 67.37 25.4 ;
        RECT 67.17 21.12 67.37 21.32 ;
        RECT 67.17 17.04 67.37 17.24 ;
        RECT 67.17 12.96 67.37 13.16 ;
        RECT 69.93 57.84 70.13 58.04 ;
        RECT 69.93 53.76 70.13 53.96 ;
        RECT 69.93 49.68 70.13 49.88 ;
        RECT 69.93 45.6 70.13 45.8 ;
        RECT 69.93 41.52 70.13 41.72 ;
        RECT 69.93 37.44 70.13 37.64 ;
        RECT 69.93 33.36 70.13 33.56 ;
        RECT 69.93 29.28 70.13 29.48 ;
        RECT 69.93 25.2 70.13 25.4 ;
        RECT 69.93 21.12 70.13 21.32 ;
        RECT 69.93 17.04 70.13 17.24 ;
        RECT 69.93 12.96 70.13 13.16 ;
        RECT 72.69 57.84 72.89 58.04 ;
        RECT 72.69 53.76 72.89 53.96 ;
        RECT 72.69 49.68 72.89 49.88 ;
        RECT 72.69 45.6 72.89 45.8 ;
        RECT 72.69 41.52 72.89 41.72 ;
        RECT 72.69 37.44 72.89 37.64 ;
        RECT 72.69 33.36 72.89 33.56 ;
        RECT 72.69 29.28 72.89 29.48 ;
        RECT 72.69 25.2 72.89 25.4 ;
        RECT 72.69 21.12 72.89 21.32 ;
        RECT 72.69 17.04 72.89 17.24 ;
        RECT 72.69 12.96 72.89 13.16 ;
        RECT 75.45 57.84 75.65 58.04 ;
        RECT 75.45 53.76 75.65 53.96 ;
        RECT 75.45 49.68 75.65 49.88 ;
        RECT 75.45 45.6 75.65 45.8 ;
        RECT 75.45 41.52 75.65 41.72 ;
        RECT 75.45 37.44 75.65 37.64 ;
        RECT 75.45 33.36 75.65 33.56 ;
        RECT 75.45 29.28 75.65 29.48 ;
        RECT 75.45 25.2 75.65 25.4 ;
        RECT 75.45 21.12 75.65 21.32 ;
        RECT 75.45 17.04 75.65 17.24 ;
        RECT 75.45 12.96 75.65 13.16 ;
        RECT 78.21 57.84 78.41 58.04 ;
        RECT 78.21 53.76 78.41 53.96 ;
        RECT 78.21 49.68 78.41 49.88 ;
        RECT 78.21 45.6 78.41 45.8 ;
        RECT 78.21 41.52 78.41 41.72 ;
        RECT 78.21 37.44 78.41 37.64 ;
        RECT 78.21 33.36 78.41 33.56 ;
        RECT 78.21 29.28 78.41 29.48 ;
        RECT 78.21 25.2 78.41 25.4 ;
        RECT 78.21 21.12 78.41 21.32 ;
        RECT 78.21 17.04 78.41 17.24 ;
        RECT 78.21 12.96 78.41 13.16 ;
        RECT 80.97 57.84 81.17 58.04 ;
        RECT 80.97 53.76 81.17 53.96 ;
        RECT 80.97 49.68 81.17 49.88 ;
        RECT 80.97 45.6 81.17 45.8 ;
        RECT 80.97 41.52 81.17 41.72 ;
        RECT 80.97 37.44 81.17 37.64 ;
        RECT 80.97 33.36 81.17 33.56 ;
        RECT 80.97 29.28 81.17 29.48 ;
        RECT 80.97 25.2 81.17 25.4 ;
        RECT 80.97 21.12 81.17 21.32 ;
        RECT 80.97 17.04 81.17 17.24 ;
        RECT 80.97 12.96 81.17 13.16 ;
        RECT 83.73 57.84 83.93 58.04 ;
        RECT 83.73 53.76 83.93 53.96 ;
        RECT 83.73 49.68 83.93 49.88 ;
        RECT 83.73 45.6 83.93 45.8 ;
        RECT 83.73 41.52 83.93 41.72 ;
        RECT 83.73 37.44 83.93 37.64 ;
        RECT 83.73 33.36 83.93 33.56 ;
        RECT 83.73 29.28 83.93 29.48 ;
        RECT 83.73 25.2 83.93 25.4 ;
        RECT 83.73 21.12 83.93 21.32 ;
        RECT 83.73 17.04 83.93 17.24 ;
        RECT 83.73 12.96 83.93 13.16 ;
        RECT 86.49 57.84 86.69 58.04 ;
        RECT 86.49 53.76 86.69 53.96 ;
        RECT 86.49 49.68 86.69 49.88 ;
        RECT 86.49 45.6 86.69 45.8 ;
        RECT 86.49 41.52 86.69 41.72 ;
        RECT 86.49 37.44 86.69 37.64 ;
        RECT 86.49 33.36 86.69 33.56 ;
        RECT 86.49 29.28 86.69 29.48 ;
        RECT 86.49 25.2 86.69 25.4 ;
        RECT 86.49 21.12 86.69 21.32 ;
        RECT 86.49 17.04 86.69 17.24 ;
        RECT 86.49 12.96 86.69 13.16 ;
        RECT 89.25 57.84 89.45 58.04 ;
        RECT 89.25 53.76 89.45 53.96 ;
        RECT 89.25 49.68 89.45 49.88 ;
        RECT 89.25 45.6 89.45 45.8 ;
        RECT 89.25 41.52 89.45 41.72 ;
        RECT 89.25 37.44 89.45 37.64 ;
        RECT 89.25 33.36 89.45 33.56 ;
        RECT 89.25 29.28 89.45 29.48 ;
        RECT 89.25 25.2 89.45 25.4 ;
        RECT 89.25 21.12 89.45 21.32 ;
        RECT 89.25 17.04 89.45 17.24 ;
        RECT 89.25 12.96 89.45 13.16 ;
        RECT 92.01 57.84 92.21 58.04 ;
        RECT 92.01 53.76 92.21 53.96 ;
        RECT 92.01 49.68 92.21 49.88 ;
        RECT 92.01 45.6 92.21 45.8 ;
        RECT 92.01 41.52 92.21 41.72 ;
        RECT 92.01 37.44 92.21 37.64 ;
        RECT 92.01 33.36 92.21 33.56 ;
        RECT 92.01 29.28 92.21 29.48 ;
        RECT 92.01 25.2 92.21 25.4 ;
        RECT 92.01 21.12 92.21 21.32 ;
        RECT 92.01 17.04 92.21 17.24 ;
        RECT 92.01 12.96 92.21 13.16 ;
        RECT 94.77 57.84 94.97 58.04 ;
        RECT 94.77 53.76 94.97 53.96 ;
        RECT 94.77 49.68 94.97 49.88 ;
        RECT 94.77 45.6 94.97 45.8 ;
        RECT 94.77 41.52 94.97 41.72 ;
        RECT 94.77 37.44 94.97 37.64 ;
        RECT 94.77 33.36 94.97 33.56 ;
        RECT 94.77 29.28 94.97 29.48 ;
        RECT 94.77 25.2 94.97 25.4 ;
        RECT 94.77 21.12 94.97 21.32 ;
        RECT 94.77 17.04 94.97 17.24 ;
        RECT 94.77 12.96 94.97 13.16 ;
        RECT 97.53 57.84 97.73 58.04 ;
        RECT 97.53 53.76 97.73 53.96 ;
        RECT 97.53 49.68 97.73 49.88 ;
        RECT 97.53 45.6 97.73 45.8 ;
        RECT 97.53 41.52 97.73 41.72 ;
        RECT 97.53 37.44 97.73 37.64 ;
        RECT 97.53 33.36 97.73 33.56 ;
        RECT 97.53 29.28 97.73 29.48 ;
        RECT 97.53 25.2 97.73 25.4 ;
        RECT 97.53 21.12 97.73 21.32 ;
        RECT 97.53 17.04 97.73 17.24 ;
        RECT 97.53 12.96 97.73 13.16 ;
        RECT 100.29 57.84 100.49 58.04 ;
        RECT 100.29 53.76 100.49 53.96 ;
        RECT 100.29 49.68 100.49 49.88 ;
        RECT 100.29 45.6 100.49 45.8 ;
        RECT 100.29 41.52 100.49 41.72 ;
        RECT 100.29 37.44 100.49 37.64 ;
        RECT 100.29 33.36 100.49 33.56 ;
        RECT 100.29 29.28 100.49 29.48 ;
        RECT 100.29 25.2 100.49 25.4 ;
        RECT 100.29 21.12 100.49 21.32 ;
        RECT 100.29 17.04 100.49 17.24 ;
        RECT 100.29 12.96 100.49 13.16 ;
        RECT 103.05 57.84 103.25 58.04 ;
        RECT 103.05 53.76 103.25 53.96 ;
        RECT 103.05 49.68 103.25 49.88 ;
        RECT 103.05 45.6 103.25 45.8 ;
        RECT 103.05 41.52 103.25 41.72 ;
        RECT 103.05 37.44 103.25 37.64 ;
        RECT 103.05 33.36 103.25 33.56 ;
        RECT 103.05 29.28 103.25 29.48 ;
        RECT 103.05 25.2 103.25 25.4 ;
        RECT 103.05 21.12 103.25 21.32 ;
        RECT 103.05 17.04 103.25 17.24 ;
        RECT 103.05 12.96 103.25 13.16 ;
        RECT 105.81 57.84 106.01 58.04 ;
        RECT 105.81 53.76 106.01 53.96 ;
        RECT 105.81 49.68 106.01 49.88 ;
        RECT 105.81 45.6 106.01 45.8 ;
        RECT 105.81 41.52 106.01 41.72 ;
        RECT 105.81 37.44 106.01 37.64 ;
        RECT 105.81 33.36 106.01 33.56 ;
        RECT 105.81 29.28 106.01 29.48 ;
        RECT 105.81 25.2 106.01 25.4 ;
        RECT 105.81 21.12 106.01 21.32 ;
        RECT 105.81 17.04 106.01 17.24 ;
        RECT 105.81 12.96 106.01 13.16 ;
        RECT 108.57 57.84 108.77 58.04 ;
        RECT 108.57 53.76 108.77 53.96 ;
        RECT 108.57 49.68 108.77 49.88 ;
        RECT 108.57 45.6 108.77 45.8 ;
        RECT 108.57 41.52 108.77 41.72 ;
        RECT 108.57 37.44 108.77 37.64 ;
        RECT 108.57 33.36 108.77 33.56 ;
        RECT 108.57 29.28 108.77 29.48 ;
        RECT 108.57 25.2 108.77 25.4 ;
        RECT 108.57 21.12 108.77 21.32 ;
        RECT 108.57 17.04 108.77 17.24 ;
        RECT 108.57 12.96 108.77 13.16 ;
        RECT 111.33 57.84 111.53 58.04 ;
        RECT 111.33 53.76 111.53 53.96 ;
        RECT 111.33 49.68 111.53 49.88 ;
        RECT 111.33 45.6 111.53 45.8 ;
        RECT 111.33 41.52 111.53 41.72 ;
        RECT 111.33 37.44 111.53 37.64 ;
        RECT 111.33 33.36 111.53 33.56 ;
        RECT 111.33 29.28 111.53 29.48 ;
        RECT 111.33 25.2 111.53 25.4 ;
        RECT 111.33 21.12 111.53 21.32 ;
        RECT 111.33 17.04 111.53 17.24 ;
        RECT 111.33 12.96 111.53 13.16 ;
        RECT 114.09 57.84 114.29 58.04 ;
        RECT 114.09 53.76 114.29 53.96 ;
        RECT 114.09 49.68 114.29 49.88 ;
        RECT 114.09 45.6 114.29 45.8 ;
        RECT 114.09 41.52 114.29 41.72 ;
        RECT 114.09 37.44 114.29 37.64 ;
        RECT 114.09 33.36 114.29 33.56 ;
        RECT 114.09 29.28 114.29 29.48 ;
        RECT 114.09 25.2 114.29 25.4 ;
        RECT 114.09 21.12 114.29 21.32 ;
        RECT 114.09 17.04 114.29 17.24 ;
        RECT 114.09 12.96 114.29 13.16 ;
        RECT 116.85 57.84 117.05 58.04 ;
        RECT 116.85 53.76 117.05 53.96 ;
        RECT 116.85 49.68 117.05 49.88 ;
        RECT 116.85 45.6 117.05 45.8 ;
        RECT 116.85 41.52 117.05 41.72 ;
        RECT 116.85 37.44 117.05 37.64 ;
        RECT 116.85 33.36 117.05 33.56 ;
        RECT 116.85 29.28 117.05 29.48 ;
        RECT 116.85 25.2 117.05 25.4 ;
        RECT 116.85 21.12 117.05 21.32 ;
        RECT 116.85 17.04 117.05 17.24 ;
        RECT 116.85 12.96 117.05 13.16 ;
        RECT 119.61 57.84 119.81 58.04 ;
        RECT 119.61 53.76 119.81 53.96 ;
        RECT 119.61 49.68 119.81 49.88 ;
        RECT 119.61 45.6 119.81 45.8 ;
        RECT 119.61 41.52 119.81 41.72 ;
        RECT 119.61 37.44 119.81 37.64 ;
        RECT 119.61 33.36 119.81 33.56 ;
        RECT 119.61 29.28 119.81 29.48 ;
        RECT 119.61 25.2 119.81 25.4 ;
        RECT 119.61 21.12 119.81 21.32 ;
        RECT 119.61 17.04 119.81 17.24 ;
        RECT 119.61 12.96 119.81 13.16 ;
        RECT 122.37 57.84 122.57 58.04 ;
        RECT 122.37 53.76 122.57 53.96 ;
        RECT 122.37 49.68 122.57 49.88 ;
        RECT 122.37 45.6 122.57 45.8 ;
        RECT 122.37 41.52 122.57 41.72 ;
        RECT 122.37 37.44 122.57 37.64 ;
        RECT 122.37 33.36 122.57 33.56 ;
        RECT 122.37 29.28 122.57 29.48 ;
        RECT 122.37 25.2 122.57 25.4 ;
        RECT 122.37 21.12 122.57 21.32 ;
        RECT 122.37 17.04 122.57 17.24 ;
        RECT 122.37 12.96 122.57 13.16 ;
        RECT 125.13 57.84 125.33 58.04 ;
        RECT 125.13 53.76 125.33 53.96 ;
        RECT 125.13 49.68 125.33 49.88 ;
        RECT 125.13 45.6 125.33 45.8 ;
        RECT 125.13 41.52 125.33 41.72 ;
        RECT 125.13 37.44 125.33 37.64 ;
        RECT 125.13 33.36 125.33 33.56 ;
        RECT 125.13 29.28 125.33 29.48 ;
        RECT 125.13 25.2 125.33 25.4 ;
        RECT 125.13 21.12 125.33 21.32 ;
        RECT 125.13 17.04 125.33 17.24 ;
        RECT 125.13 12.96 125.33 13.16 ;
        RECT 127.89 57.84 128.09 58.04 ;
        RECT 127.89 53.76 128.09 53.96 ;
        RECT 127.89 49.68 128.09 49.88 ;
        RECT 127.89 45.6 128.09 45.8 ;
        RECT 127.89 41.52 128.09 41.72 ;
        RECT 127.89 37.44 128.09 37.64 ;
        RECT 127.89 33.36 128.09 33.56 ;
        RECT 127.89 29.28 128.09 29.48 ;
        RECT 127.89 25.2 128.09 25.4 ;
        RECT 127.89 21.12 128.09 21.32 ;
        RECT 127.89 17.04 128.09 17.24 ;
        RECT 127.89 12.96 128.09 13.16 ;
        RECT 130.65 57.84 130.85 58.04 ;
        RECT 130.65 53.76 130.85 53.96 ;
        RECT 130.65 49.68 130.85 49.88 ;
        RECT 130.65 45.6 130.85 45.8 ;
        RECT 130.65 41.52 130.85 41.72 ;
        RECT 130.65 37.44 130.85 37.64 ;
        RECT 130.65 33.36 130.85 33.56 ;
        RECT 130.65 29.28 130.85 29.48 ;
        RECT 130.65 25.2 130.85 25.4 ;
        RECT 130.65 21.12 130.85 21.32 ;
        RECT 130.65 17.04 130.85 17.24 ;
        RECT 130.65 12.96 130.85 13.16 ;
        RECT 133.41 57.84 133.61 58.04 ;
        RECT 133.41 53.76 133.61 53.96 ;
        RECT 133.41 49.68 133.61 49.88 ;
        RECT 133.41 45.6 133.61 45.8 ;
        RECT 133.41 41.52 133.61 41.72 ;
        RECT 133.41 37.44 133.61 37.64 ;
        RECT 133.41 33.36 133.61 33.56 ;
        RECT 133.41 29.28 133.61 29.48 ;
        RECT 133.41 25.2 133.61 25.4 ;
        RECT 133.41 21.12 133.61 21.32 ;
        RECT 133.41 17.04 133.61 17.24 ;
        RECT 133.41 12.96 133.61 13.16 ;
        RECT 136.17 57.84 136.37 58.04 ;
        RECT 136.17 53.76 136.37 53.96 ;
        RECT 136.17 49.68 136.37 49.88 ;
        RECT 136.17 45.6 136.37 45.8 ;
        RECT 136.17 41.52 136.37 41.72 ;
        RECT 136.17 37.44 136.37 37.64 ;
        RECT 136.17 33.36 136.37 33.56 ;
        RECT 136.17 29.28 136.37 29.48 ;
        RECT 136.17 25.2 136.37 25.4 ;
        RECT 136.17 21.12 136.37 21.32 ;
        RECT 136.17 17.04 136.37 17.24 ;
        RECT 136.17 12.96 136.37 13.16 ;
        RECT 138.93 57.84 139.13 58.04 ;
        RECT 138.93 53.76 139.13 53.96 ;
        RECT 138.93 49.68 139.13 49.88 ;
        RECT 138.93 45.6 139.13 45.8 ;
        RECT 138.93 41.52 139.13 41.72 ;
        RECT 138.93 37.44 139.13 37.64 ;
        RECT 138.93 33.36 139.13 33.56 ;
        RECT 138.93 29.28 139.13 29.48 ;
        RECT 138.93 25.2 139.13 25.4 ;
        RECT 138.93 21.12 139.13 21.32 ;
        RECT 138.93 17.04 139.13 17.24 ;
        RECT 138.93 12.96 139.13 13.16 ;
        RECT 141.69 57.84 141.89 58.04 ;
        RECT 141.69 53.76 141.89 53.96 ;
        RECT 141.69 49.68 141.89 49.88 ;
        RECT 141.69 45.6 141.89 45.8 ;
        RECT 141.69 41.52 141.89 41.72 ;
        RECT 141.69 37.44 141.89 37.64 ;
        RECT 141.69 33.36 141.89 33.56 ;
        RECT 141.69 29.28 141.89 29.48 ;
        RECT 141.69 25.2 141.89 25.4 ;
        RECT 141.69 21.12 141.89 21.32 ;
        RECT 141.69 17.04 141.89 17.24 ;
        RECT 141.69 12.96 141.89 13.16 ;
        RECT 144.45 57.84 144.65 58.04 ;
        RECT 144.45 53.76 144.65 53.96 ;
        RECT 144.45 49.68 144.65 49.88 ;
        RECT 144.45 45.6 144.65 45.8 ;
        RECT 144.45 41.52 144.65 41.72 ;
        RECT 144.45 37.44 144.65 37.64 ;
        RECT 144.45 33.36 144.65 33.56 ;
        RECT 144.45 29.28 144.65 29.48 ;
        RECT 144.45 25.2 144.65 25.4 ;
        RECT 144.45 21.12 144.65 21.32 ;
        RECT 144.45 17.04 144.65 17.24 ;
        RECT 144.45 12.96 144.65 13.16 ;
        RECT 147.21 57.84 147.41 58.04 ;
        RECT 147.21 53.76 147.41 53.96 ;
        RECT 147.21 49.68 147.41 49.88 ;
        RECT 147.21 45.6 147.41 45.8 ;
        RECT 147.21 41.52 147.41 41.72 ;
        RECT 147.21 37.44 147.41 37.64 ;
        RECT 147.21 33.36 147.41 33.56 ;
        RECT 147.21 29.28 147.41 29.48 ;
        RECT 147.21 25.2 147.41 25.4 ;
        RECT 147.21 21.12 147.41 21.32 ;
        RECT 147.21 17.04 147.41 17.24 ;
        RECT 147.21 12.96 147.41 13.16 ;
        RECT 149.97 57.84 150.17 58.04 ;
        RECT 149.97 53.76 150.17 53.96 ;
        RECT 149.97 49.68 150.17 49.88 ;
        RECT 149.97 45.6 150.17 45.8 ;
        RECT 149.97 41.52 150.17 41.72 ;
        RECT 149.97 37.44 150.17 37.64 ;
        RECT 149.97 33.36 150.17 33.56 ;
        RECT 149.97 29.28 150.17 29.48 ;
        RECT 149.97 25.2 150.17 25.4 ;
        RECT 149.97 21.12 150.17 21.32 ;
        RECT 149.97 17.04 150.17 17.24 ;
        RECT 149.97 12.96 150.17 13.16 ;
        RECT 152.73 57.84 152.93 58.04 ;
        RECT 152.73 53.76 152.93 53.96 ;
        RECT 152.73 49.68 152.93 49.88 ;
        RECT 152.73 45.6 152.93 45.8 ;
        RECT 152.73 41.52 152.93 41.72 ;
        RECT 152.73 37.44 152.93 37.64 ;
        RECT 152.73 33.36 152.93 33.56 ;
        RECT 152.73 29.28 152.93 29.48 ;
        RECT 152.73 25.2 152.93 25.4 ;
        RECT 152.73 21.12 152.93 21.32 ;
        RECT 152.73 17.04 152.93 17.24 ;
        RECT 152.73 12.96 152.93 13.16 ;
        RECT 155.49 57.84 155.69 58.04 ;
        RECT 155.49 53.76 155.69 53.96 ;
        RECT 155.49 49.68 155.69 49.88 ;
        RECT 155.49 45.6 155.69 45.8 ;
        RECT 155.49 41.52 155.69 41.72 ;
        RECT 155.49 37.44 155.69 37.64 ;
        RECT 155.49 33.36 155.69 33.56 ;
        RECT 155.49 29.28 155.69 29.48 ;
        RECT 155.49 25.2 155.69 25.4 ;
        RECT 155.49 21.12 155.69 21.32 ;
        RECT 155.49 17.04 155.69 17.24 ;
        RECT 155.49 12.96 155.69 13.16 ;
        RECT 158.25 57.84 158.45 58.04 ;
        RECT 158.25 53.76 158.45 53.96 ;
        RECT 158.25 49.68 158.45 49.88 ;
        RECT 158.25 45.6 158.45 45.8 ;
        RECT 158.25 41.52 158.45 41.72 ;
        RECT 158.25 37.44 158.45 37.64 ;
        RECT 158.25 33.36 158.45 33.56 ;
        RECT 158.25 29.28 158.45 29.48 ;
        RECT 158.25 25.2 158.45 25.4 ;
        RECT 158.25 21.12 158.45 21.32 ;
        RECT 158.25 17.04 158.45 17.24 ;
        RECT 158.25 12.96 158.45 13.16 ;
        RECT 161.01 57.84 161.21 58.04 ;
        RECT 161.01 53.76 161.21 53.96 ;
        RECT 161.01 49.68 161.21 49.88 ;
        RECT 161.01 45.6 161.21 45.8 ;
        RECT 161.01 41.52 161.21 41.72 ;
        RECT 161.01 37.44 161.21 37.64 ;
        RECT 161.01 33.36 161.21 33.56 ;
        RECT 161.01 29.28 161.21 29.48 ;
        RECT 161.01 25.2 161.21 25.4 ;
        RECT 161.01 21.12 161.21 21.32 ;
        RECT 161.01 17.04 161.21 17.24 ;
        RECT 161.01 12.96 161.21 13.16 ;
        RECT 163.77 57.84 163.97 58.04 ;
        RECT 163.77 53.76 163.97 53.96 ;
        RECT 163.77 49.68 163.97 49.88 ;
        RECT 163.77 45.6 163.97 45.8 ;
        RECT 163.77 41.52 163.97 41.72 ;
        RECT 163.77 37.44 163.97 37.64 ;
        RECT 163.77 33.36 163.97 33.56 ;
        RECT 163.77 29.28 163.97 29.48 ;
        RECT 163.77 25.2 163.97 25.4 ;
        RECT 163.77 21.12 163.97 21.32 ;
        RECT 163.77 17.04 163.97 17.24 ;
        RECT 163.77 12.96 163.97 13.16 ;
        RECT 166.53 57.84 166.73 58.04 ;
        RECT 166.53 53.76 166.73 53.96 ;
        RECT 166.53 49.68 166.73 49.88 ;
        RECT 166.53 45.6 166.73 45.8 ;
        RECT 166.53 41.52 166.73 41.72 ;
        RECT 166.53 37.44 166.73 37.64 ;
        RECT 166.53 33.36 166.73 33.56 ;
        RECT 166.53 29.28 166.73 29.48 ;
        RECT 166.53 25.2 166.73 25.4 ;
        RECT 166.53 21.12 166.73 21.32 ;
        RECT 166.53 17.04 166.73 17.24 ;
        RECT 166.53 12.96 166.73 13.16 ;
        RECT 169.29 57.84 169.49 58.04 ;
        RECT 169.29 53.76 169.49 53.96 ;
        RECT 169.29 49.68 169.49 49.88 ;
        RECT 169.29 45.6 169.49 45.8 ;
        RECT 169.29 41.52 169.49 41.72 ;
        RECT 169.29 37.44 169.49 37.64 ;
        RECT 169.29 33.36 169.49 33.56 ;
        RECT 169.29 29.28 169.49 29.48 ;
        RECT 169.29 25.2 169.49 25.4 ;
        RECT 169.29 21.12 169.49 21.32 ;
        RECT 169.29 17.04 169.49 17.24 ;
        RECT 169.29 12.96 169.49 13.16 ;
        RECT 172.05 57.84 172.25 58.04 ;
        RECT 172.05 53.76 172.25 53.96 ;
        RECT 172.05 49.68 172.25 49.88 ;
        RECT 172.05 45.6 172.25 45.8 ;
        RECT 172.05 41.52 172.25 41.72 ;
        RECT 172.05 37.44 172.25 37.64 ;
        RECT 172.05 33.36 172.25 33.56 ;
        RECT 172.05 29.28 172.25 29.48 ;
        RECT 172.05 25.2 172.25 25.4 ;
        RECT 172.05 21.12 172.25 21.32 ;
        RECT 172.05 17.04 172.25 17.24 ;
        RECT 172.05 12.96 172.25 13.16 ;
        RECT 174.81 57.84 175.01 58.04 ;
        RECT 174.81 53.76 175.01 53.96 ;
        RECT 174.81 49.68 175.01 49.88 ;
        RECT 174.81 45.6 175.01 45.8 ;
        RECT 174.81 41.52 175.01 41.72 ;
        RECT 174.81 37.44 175.01 37.64 ;
        RECT 174.81 33.36 175.01 33.56 ;
        RECT 174.81 29.28 175.01 29.48 ;
        RECT 174.81 25.2 175.01 25.4 ;
        RECT 174.81 21.12 175.01 21.32 ;
        RECT 174.81 17.04 175.01 17.24 ;
        RECT 174.81 12.96 175.01 13.16 ;
        RECT 177.57 57.84 177.77 58.04 ;
        RECT 177.57 53.76 177.77 53.96 ;
        RECT 177.57 49.68 177.77 49.88 ;
        RECT 177.57 45.6 177.77 45.8 ;
        RECT 177.57 41.52 177.77 41.72 ;
        RECT 177.57 37.44 177.77 37.64 ;
        RECT 177.57 33.36 177.77 33.56 ;
        RECT 177.57 29.28 177.77 29.48 ;
        RECT 177.57 25.2 177.77 25.4 ;
        RECT 177.57 21.12 177.77 21.32 ;
        RECT 177.57 17.04 177.77 17.24 ;
        RECT 177.57 12.96 177.77 13.16 ;
        RECT 180.33 57.84 180.53 58.04 ;
        RECT 180.33 53.76 180.53 53.96 ;
        RECT 180.33 49.68 180.53 49.88 ;
        RECT 180.33 45.6 180.53 45.8 ;
        RECT 180.33 41.52 180.53 41.72 ;
        RECT 180.33 37.44 180.53 37.64 ;
        RECT 180.33 33.36 180.53 33.56 ;
        RECT 180.33 29.28 180.53 29.48 ;
        RECT 180.33 25.2 180.53 25.4 ;
        RECT 180.33 21.12 180.53 21.32 ;
        RECT 180.33 17.04 180.53 17.24 ;
        RECT 180.33 12.96 180.53 13.16 ;
        RECT 183.09 57.84 183.29 58.04 ;
        RECT 183.09 53.76 183.29 53.96 ;
        RECT 183.09 49.68 183.29 49.88 ;
        RECT 183.09 45.6 183.29 45.8 ;
        RECT 183.09 41.52 183.29 41.72 ;
        RECT 183.09 37.44 183.29 37.64 ;
        RECT 183.09 33.36 183.29 33.56 ;
        RECT 183.09 29.28 183.29 29.48 ;
        RECT 183.09 25.2 183.29 25.4 ;
        RECT 183.09 21.12 183.29 21.32 ;
        RECT 183.09 17.04 183.29 17.24 ;
        RECT 183.09 12.96 183.29 13.16 ;
        RECT 185.85 57.84 186.05 58.04 ;
        RECT 185.85 53.76 186.05 53.96 ;
        RECT 185.85 49.68 186.05 49.88 ;
        RECT 185.85 45.6 186.05 45.8 ;
        RECT 185.85 41.52 186.05 41.72 ;
        RECT 185.85 37.44 186.05 37.64 ;
        RECT 185.85 33.36 186.05 33.56 ;
        RECT 185.85 29.28 186.05 29.48 ;
        RECT 185.85 25.2 186.05 25.4 ;
        RECT 185.85 21.12 186.05 21.32 ;
        RECT 185.85 17.04 186.05 17.24 ;
        RECT 185.85 12.96 186.05 13.16 ;
        RECT 188.61 57.84 188.81 58.04 ;
        RECT 188.61 53.76 188.81 53.96 ;
        RECT 188.61 49.68 188.81 49.88 ;
        RECT 188.61 45.6 188.81 45.8 ;
        RECT 188.61 41.52 188.81 41.72 ;
        RECT 188.61 37.44 188.81 37.64 ;
        RECT 188.61 33.36 188.81 33.56 ;
        RECT 188.61 29.28 188.81 29.48 ;
        RECT 188.61 25.2 188.81 25.4 ;
        RECT 188.61 21.12 188.81 21.32 ;
        RECT 188.61 17.04 188.81 17.24 ;
        RECT 188.61 12.96 188.81 13.16 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met5 ;
        RECT 0 17.5 200 19.5 ;
        RECT 0 37.9 200 39.9 ;
      LAYER li1 ;
        RECT 79.545 33.625 84.89 35.335 ;
        RECT 79.545 33.105 82.125 35.855 ;
        RECT 74.025 33.625 79.37 35.335 ;
        RECT 74.025 33.105 76.605 35.855 ;
        RECT 73.565 33.67 73.855 35.29 ;
        RECT 72.185 33.645 73.395 35.315 ;
        RECT 72.185 33.105 72.705 35.855 ;
        RECT 70.345 33.625 72.015 35.335 ;
        RECT 70.345 33.105 71.095 35.855 ;
        RECT 64.825 33.625 70.17 35.335 ;
        RECT 64.825 33.105 67.405 35.855 ;
        RECT 59.305 33.625 64.65 35.335 ;
        RECT 59.305 33.105 61.885 35.855 ;
        RECT 58.845 33.67 59.135 35.29 ;
        RECT 57.465 33.625 58.675 35.315 ;
        RECT 57.465 33.625 57.985 35.855 ;
        RECT 56.085 33.625 58.675 34.565 ;
        RECT 56.085 33.105 57.295 35.335 ;
        RECT 55.625 34.395 56.375 35.855 ;
        RECT 55.195 33.785 55.365 34.565 ;
        RECT 54.735 34.395 54.905 35.175 ;
        RECT 54.225 33.865 54.435 34.565 ;
        RECT 53.765 34.395 53.975 35.095 ;
        RECT 52.04 33.895 52.41 34.565 ;
        RECT 51.58 34.395 51.95 35.065 ;
        RECT 50.095 33.935 50.345 34.565 ;
        RECT 49.635 34.395 49.885 35.025 ;
        RECT 49.155 34.015 49.485 34.565 ;
        RECT 48.695 34.395 49.025 34.945 ;
        RECT 47.345 33.645 48.555 34.565 ;
        RECT 44.585 34.395 48.095 35.335 ;
        RECT 47.345 33.105 47.865 35.335 ;
        RECT 44.585 33.625 47.175 35.335 ;
        RECT 44.585 33.625 46.235 35.855 ;
        RECT 44.585 33.105 45.795 35.855 ;
        RECT 44.125 33.67 44.415 35.29 ;
        RECT 42.745 33.645 43.955 35.315 ;
        RECT 42.745 33.105 43.265 35.855 ;
        RECT 40.905 33.625 42.575 35.335 ;
        RECT 40.905 33.105 41.655 35.855 ;
        RECT 35.385 33.625 40.73 35.335 ;
        RECT 35.385 33.105 37.965 35.855 ;
        RECT 29.865 33.625 35.21 35.335 ;
        RECT 29.865 33.105 32.445 35.855 ;
        RECT 29.405 33.67 29.695 35.29 ;
        RECT 28.025 33.645 29.235 35.315 ;
        RECT 28.025 33.105 28.545 35.855 ;
        RECT 26.185 33.625 27.855 35.335 ;
        RECT 26.185 33.105 26.935 35.855 ;
        RECT 20.665 33.625 26.01 35.335 ;
        RECT 20.665 33.105 23.245 35.855 ;
        RECT 15.145 33.625 20.49 35.335 ;
        RECT 15.145 33.105 17.725 35.855 ;
        RECT 14.685 33.67 14.975 35.29 ;
        RECT 13.305 33.645 14.515 35.315 ;
        RECT 13.305 33.105 13.825 35.855 ;
        RECT 10.545 33.625 13.135 35.335 ;
        RECT 10.545 33.105 11.755 35.855 ;
        RECT 10 39.835 189.86 40.005 ;
        RECT 189.025 39.11 189.315 40.73 ;
        RECT 186.265 39.065 188.855 40.775 ;
        RECT 186.265 38.545 187.475 41.295 ;
        RECT 182.585 39.065 186.095 40.775 ;
        RECT 182.585 38.545 184.235 41.295 ;
        RECT 177.065 39.065 182.41 40.775 ;
        RECT 177.065 38.545 179.645 41.295 ;
        RECT 176.605 39.11 176.895 40.73 ;
        RECT 175.225 39.085 176.435 40.755 ;
        RECT 175.225 38.545 175.745 41.295 ;
        RECT 173.385 39.065 175.055 40.775 ;
        RECT 173.385 38.545 174.135 41.295 ;
        RECT 167.865 39.065 173.21 40.775 ;
        RECT 167.865 38.545 170.445 41.295 ;
        RECT 162.345 39.065 167.69 40.775 ;
        RECT 162.345 38.545 164.925 41.295 ;
        RECT 161.885 39.11 162.175 40.73 ;
        RECT 160.505 39.085 161.715 40.755 ;
        RECT 160.505 38.545 161.025 41.295 ;
        RECT 158.665 39.065 160.335 40.775 ;
        RECT 158.665 38.545 159.415 41.295 ;
        RECT 153.145 39.065 158.49 40.775 ;
        RECT 153.145 38.545 155.725 41.295 ;
        RECT 147.625 39.065 152.97 40.775 ;
        RECT 147.625 38.545 150.205 41.295 ;
        RECT 147.165 39.11 147.455 40.73 ;
        RECT 145.785 39.085 146.995 40.755 ;
        RECT 145.785 38.545 146.305 41.295 ;
        RECT 143.945 39.065 145.615 40.775 ;
        RECT 143.945 38.545 144.695 41.295 ;
        RECT 138.425 39.065 143.77 40.775 ;
        RECT 138.425 38.545 141.005 41.295 ;
        RECT 132.905 39.065 138.25 40.775 ;
        RECT 132.905 38.545 135.485 41.295 ;
        RECT 132.445 39.11 132.735 40.73 ;
        RECT 131.065 39.085 132.275 40.755 ;
        RECT 131.065 38.545 131.585 41.295 ;
        RECT 129.225 39.065 130.895 40.775 ;
        RECT 129.225 38.545 129.975 41.295 ;
        RECT 123.705 39.065 129.05 40.775 ;
        RECT 123.705 38.545 126.285 41.295 ;
        RECT 118.185 39.065 123.53 40.775 ;
        RECT 118.185 38.545 120.765 41.295 ;
        RECT 117.725 39.11 118.015 40.73 ;
        RECT 116.345 39.085 117.555 40.755 ;
        RECT 116.345 38.545 116.865 41.295 ;
        RECT 114.505 39.065 116.175 40.775 ;
        RECT 114.505 38.545 115.255 41.295 ;
        RECT 108.985 39.065 114.33 40.775 ;
        RECT 108.985 38.545 111.565 41.295 ;
        RECT 103.465 39.065 108.81 40.775 ;
        RECT 103.465 38.545 106.045 41.295 ;
        RECT 103.005 39.11 103.295 40.73 ;
        RECT 101.625 39.085 102.835 40.755 ;
        RECT 101.625 38.545 102.145 41.295 ;
        RECT 99.785 39.065 101.455 40.775 ;
        RECT 99.785 38.545 100.535 41.295 ;
        RECT 94.265 39.065 99.61 40.775 ;
        RECT 94.265 38.545 96.845 41.295 ;
        RECT 88.745 39.065 94.09 40.775 ;
        RECT 88.745 38.545 91.325 41.295 ;
        RECT 88.285 39.11 88.575 40.73 ;
        RECT 86.905 39.085 88.115 40.755 ;
        RECT 86.905 38.545 87.425 41.295 ;
        RECT 85.065 39.065 86.735 40.775 ;
        RECT 85.065 38.545 85.815 41.295 ;
        RECT 79.545 39.065 84.89 40.775 ;
        RECT 79.545 38.545 82.125 41.295 ;
        RECT 74.025 39.065 79.37 40.775 ;
        RECT 74.025 38.545 76.605 41.295 ;
        RECT 73.565 39.11 73.855 40.73 ;
        RECT 72.185 39.085 73.395 40.755 ;
        RECT 72.185 38.545 72.705 41.295 ;
        RECT 70.345 39.065 72.015 40.775 ;
        RECT 70.345 38.545 71.095 41.295 ;
        RECT 64.825 39.065 70.17 40.775 ;
        RECT 64.825 38.545 67.405 41.295 ;
        RECT 59.305 39.065 64.65 40.775 ;
        RECT 59.305 38.545 61.885 41.295 ;
        RECT 58.845 39.11 59.135 40.73 ;
        RECT 57.465 39.085 58.675 40.755 ;
        RECT 57.465 38.545 57.985 41.295 ;
        RECT 55.625 39.065 57.295 40.775 ;
        RECT 55.625 38.545 56.375 41.295 ;
        RECT 50.105 39.065 55.45 40.775 ;
        RECT 50.105 38.545 52.685 41.295 ;
        RECT 44.585 39.065 49.93 40.775 ;
        RECT 44.585 38.545 47.165 41.295 ;
        RECT 44.125 39.11 44.415 40.73 ;
        RECT 42.745 39.085 43.955 40.755 ;
        RECT 42.745 38.545 43.265 41.295 ;
        RECT 40.905 39.065 42.575 40.775 ;
        RECT 40.905 38.545 41.655 41.295 ;
        RECT 35.385 39.065 40.73 40.775 ;
        RECT 35.385 38.545 37.965 41.295 ;
        RECT 29.865 39.065 35.21 40.775 ;
        RECT 29.865 38.545 32.445 41.295 ;
        RECT 29.405 39.11 29.695 40.73 ;
        RECT 28.025 39.085 29.235 40.755 ;
        RECT 28.025 38.545 28.545 41.295 ;
        RECT 26.185 39.065 27.855 40.775 ;
        RECT 26.185 38.545 26.935 41.295 ;
        RECT 20.665 39.065 26.01 40.775 ;
        RECT 20.665 38.545 23.245 41.295 ;
        RECT 15.145 39.065 20.49 40.775 ;
        RECT 15.145 38.545 17.725 41.295 ;
        RECT 14.685 39.11 14.975 40.73 ;
        RECT 13.305 39.085 14.515 40.755 ;
        RECT 13.305 38.545 13.825 41.295 ;
        RECT 10.545 39.065 13.135 40.775 ;
        RECT 10.545 38.545 11.755 41.295 ;
        RECT 10 45.275 189.86 45.445 ;
        RECT 189.025 44.55 189.315 46.17 ;
        RECT 186.265 44.505 188.855 46.215 ;
        RECT 186.265 43.985 187.475 46.735 ;
        RECT 182.585 44.505 186.095 46.215 ;
        RECT 182.585 43.985 184.235 46.735 ;
        RECT 177.065 44.505 182.41 46.215 ;
        RECT 177.065 43.985 179.645 46.735 ;
        RECT 176.605 44.55 176.895 46.17 ;
        RECT 175.225 44.525 176.435 46.195 ;
        RECT 175.225 43.985 175.745 46.735 ;
        RECT 173.385 44.505 175.055 46.215 ;
        RECT 173.385 43.985 174.135 46.735 ;
        RECT 167.865 44.505 173.21 46.215 ;
        RECT 167.865 43.985 170.445 46.735 ;
        RECT 162.345 44.505 167.69 46.215 ;
        RECT 162.345 43.985 164.925 46.735 ;
        RECT 161.885 44.55 162.175 46.17 ;
        RECT 160.505 44.525 161.715 46.195 ;
        RECT 160.505 43.985 161.025 46.735 ;
        RECT 158.665 44.505 160.335 46.215 ;
        RECT 158.665 43.985 159.415 46.735 ;
        RECT 153.145 44.505 158.49 46.215 ;
        RECT 153.145 43.985 155.725 46.735 ;
        RECT 147.625 44.505 152.97 46.215 ;
        RECT 147.625 43.985 150.205 46.735 ;
        RECT 147.165 44.55 147.455 46.17 ;
        RECT 145.785 44.525 146.995 46.195 ;
        RECT 145.785 43.985 146.305 46.735 ;
        RECT 143.945 44.505 145.615 46.215 ;
        RECT 143.945 43.985 144.695 46.735 ;
        RECT 138.425 44.505 143.77 46.215 ;
        RECT 138.425 43.985 141.005 46.735 ;
        RECT 132.905 44.505 138.25 46.215 ;
        RECT 132.905 43.985 135.485 46.735 ;
        RECT 132.445 44.55 132.735 46.17 ;
        RECT 131.065 44.525 132.275 46.195 ;
        RECT 131.065 43.985 131.585 46.735 ;
        RECT 129.225 44.505 130.895 46.215 ;
        RECT 129.225 43.985 129.975 46.735 ;
        RECT 123.705 44.505 129.05 46.215 ;
        RECT 123.705 43.985 126.285 46.735 ;
        RECT 118.185 44.505 123.53 46.215 ;
        RECT 118.185 43.985 120.765 46.735 ;
        RECT 117.725 44.55 118.015 46.17 ;
        RECT 116.345 44.525 117.555 46.195 ;
        RECT 116.345 43.985 116.865 46.735 ;
        RECT 114.505 44.505 116.175 46.215 ;
        RECT 114.505 43.985 115.255 46.735 ;
        RECT 108.985 44.505 114.33 46.215 ;
        RECT 108.985 43.985 111.565 46.735 ;
        RECT 103.465 44.505 108.81 46.215 ;
        RECT 103.465 43.985 106.045 46.735 ;
        RECT 103.005 44.55 103.295 46.17 ;
        RECT 101.625 44.525 102.835 46.195 ;
        RECT 101.625 43.985 102.145 46.735 ;
        RECT 99.785 44.505 101.455 46.215 ;
        RECT 99.785 43.985 100.535 46.735 ;
        RECT 94.265 44.505 99.61 46.215 ;
        RECT 94.265 43.985 96.845 46.735 ;
        RECT 88.745 44.505 94.09 46.215 ;
        RECT 88.745 43.985 91.325 46.735 ;
        RECT 88.285 44.55 88.575 46.17 ;
        RECT 86.905 44.525 88.115 46.195 ;
        RECT 86.905 43.985 87.425 46.735 ;
        RECT 85.065 44.505 86.735 46.215 ;
        RECT 85.065 43.985 85.815 46.735 ;
        RECT 79.545 44.505 84.89 46.215 ;
        RECT 79.545 43.985 82.125 46.735 ;
        RECT 74.025 44.505 79.37 46.215 ;
        RECT 74.025 43.985 76.605 46.735 ;
        RECT 73.565 44.55 73.855 46.17 ;
        RECT 72.185 44.525 73.395 46.195 ;
        RECT 72.185 43.985 72.705 46.735 ;
        RECT 70.345 44.505 72.015 46.215 ;
        RECT 70.345 43.985 71.095 46.735 ;
        RECT 64.825 44.505 70.17 46.215 ;
        RECT 64.825 43.985 67.405 46.735 ;
        RECT 59.305 44.505 64.65 46.215 ;
        RECT 59.305 43.985 61.885 46.735 ;
        RECT 58.845 44.55 59.135 46.17 ;
        RECT 57.465 44.525 58.675 46.195 ;
        RECT 57.465 43.985 57.985 46.735 ;
        RECT 55.625 44.505 57.295 46.215 ;
        RECT 55.625 43.985 56.375 46.735 ;
        RECT 50.105 44.505 55.45 46.215 ;
        RECT 50.105 43.985 52.685 46.735 ;
        RECT 44.585 44.505 49.93 46.215 ;
        RECT 44.585 43.985 47.165 46.735 ;
        RECT 44.125 44.55 44.415 46.17 ;
        RECT 42.745 44.525 43.955 46.195 ;
        RECT 42.745 43.985 43.265 46.735 ;
        RECT 40.905 44.505 42.575 46.215 ;
        RECT 40.905 43.985 41.655 46.735 ;
        RECT 35.385 44.505 40.73 46.215 ;
        RECT 35.385 43.985 37.965 46.735 ;
        RECT 29.865 44.505 35.21 46.215 ;
        RECT 29.865 43.985 32.445 46.735 ;
        RECT 29.405 44.55 29.695 46.17 ;
        RECT 28.025 44.525 29.235 46.195 ;
        RECT 28.025 43.985 28.545 46.735 ;
        RECT 26.185 44.505 27.855 46.215 ;
        RECT 26.185 43.985 26.935 46.735 ;
        RECT 20.665 44.505 26.01 46.215 ;
        RECT 20.665 43.985 23.245 46.735 ;
        RECT 15.145 44.505 20.49 46.215 ;
        RECT 15.145 43.985 17.725 46.735 ;
        RECT 14.685 44.55 14.975 46.17 ;
        RECT 13.305 44.525 14.515 46.195 ;
        RECT 13.305 43.985 13.825 46.735 ;
        RECT 10.545 44.505 13.135 46.215 ;
        RECT 10.545 43.985 11.755 46.735 ;
        RECT 10 50.715 189.86 50.885 ;
        RECT 189.025 49.99 189.315 51.61 ;
        RECT 186.265 49.945 188.855 51.655 ;
        RECT 186.265 49.425 187.475 52.175 ;
        RECT 182.585 49.945 186.095 51.655 ;
        RECT 182.585 49.425 184.235 52.175 ;
        RECT 177.065 49.945 182.41 51.655 ;
        RECT 177.065 49.425 179.645 52.175 ;
        RECT 176.605 49.99 176.895 51.61 ;
        RECT 175.225 49.965 176.435 51.635 ;
        RECT 175.225 49.425 175.745 52.175 ;
        RECT 173.385 49.945 175.055 51.655 ;
        RECT 173.385 49.425 174.135 52.175 ;
        RECT 167.865 49.945 173.21 51.655 ;
        RECT 167.865 49.425 170.445 52.175 ;
        RECT 162.345 49.945 167.69 51.655 ;
        RECT 162.345 49.425 164.925 52.175 ;
        RECT 161.885 49.99 162.175 51.61 ;
        RECT 160.505 49.965 161.715 51.635 ;
        RECT 160.505 49.425 161.025 52.175 ;
        RECT 158.665 49.945 160.335 51.655 ;
        RECT 158.665 49.425 159.415 52.175 ;
        RECT 153.145 49.945 158.49 51.655 ;
        RECT 153.145 49.425 155.725 52.175 ;
        RECT 147.625 49.945 152.97 51.655 ;
        RECT 147.625 49.425 150.205 52.175 ;
        RECT 147.165 49.99 147.455 51.61 ;
        RECT 145.785 49.965 146.995 51.635 ;
        RECT 145.785 49.425 146.305 52.175 ;
        RECT 143.945 49.945 145.615 51.655 ;
        RECT 143.945 49.425 144.695 52.175 ;
        RECT 138.425 49.945 143.77 51.655 ;
        RECT 138.425 49.425 141.005 52.175 ;
        RECT 132.905 49.945 138.25 51.655 ;
        RECT 132.905 49.425 135.485 52.175 ;
        RECT 132.445 49.99 132.735 51.61 ;
        RECT 131.065 49.965 132.275 51.635 ;
        RECT 131.065 49.425 131.585 52.175 ;
        RECT 129.225 49.945 130.895 51.655 ;
        RECT 129.225 49.425 129.975 52.175 ;
        RECT 123.705 49.945 129.05 51.655 ;
        RECT 123.705 49.425 126.285 52.175 ;
        RECT 118.185 49.945 123.53 51.655 ;
        RECT 118.185 49.425 120.765 52.175 ;
        RECT 117.725 49.99 118.015 51.61 ;
        RECT 116.345 49.965 117.555 51.635 ;
        RECT 116.345 49.425 116.865 52.175 ;
        RECT 114.505 49.945 116.175 51.655 ;
        RECT 114.505 49.425 115.255 52.175 ;
        RECT 108.985 49.945 114.33 51.655 ;
        RECT 108.985 49.425 111.565 52.175 ;
        RECT 103.465 49.945 108.81 51.655 ;
        RECT 103.465 49.425 106.045 52.175 ;
        RECT 103.005 49.99 103.295 51.61 ;
        RECT 101.625 49.965 102.835 51.635 ;
        RECT 101.625 49.425 102.145 52.175 ;
        RECT 99.785 49.945 101.455 51.655 ;
        RECT 99.785 49.425 100.535 52.175 ;
        RECT 94.265 49.945 99.61 51.655 ;
        RECT 94.265 49.425 96.845 52.175 ;
        RECT 88.745 49.945 94.09 51.655 ;
        RECT 88.745 49.425 91.325 52.175 ;
        RECT 88.285 49.99 88.575 51.61 ;
        RECT 86.905 49.965 88.115 51.635 ;
        RECT 86.905 49.425 87.425 52.175 ;
        RECT 85.065 49.945 86.735 51.655 ;
        RECT 85.065 49.425 85.815 52.175 ;
        RECT 79.545 49.945 84.89 51.655 ;
        RECT 79.545 49.425 82.125 52.175 ;
        RECT 74.025 49.945 79.37 51.655 ;
        RECT 74.025 49.425 76.605 52.175 ;
        RECT 73.565 49.99 73.855 51.61 ;
        RECT 72.185 49.965 73.395 51.635 ;
        RECT 72.185 49.425 72.705 52.175 ;
        RECT 70.345 49.945 72.015 51.655 ;
        RECT 70.345 49.425 71.095 52.175 ;
        RECT 64.825 49.945 70.17 51.655 ;
        RECT 64.825 49.425 67.405 52.175 ;
        RECT 59.305 49.945 64.65 51.655 ;
        RECT 59.305 49.425 61.885 52.175 ;
        RECT 58.845 49.99 59.135 51.61 ;
        RECT 57.465 49.965 58.675 51.635 ;
        RECT 57.465 49.425 57.985 52.175 ;
        RECT 55.625 49.945 57.295 51.655 ;
        RECT 55.625 49.425 56.375 52.175 ;
        RECT 50.105 49.945 55.45 51.655 ;
        RECT 50.105 49.425 52.685 52.175 ;
        RECT 44.585 49.945 49.93 51.655 ;
        RECT 44.585 49.425 47.165 52.175 ;
        RECT 44.125 49.99 44.415 51.61 ;
        RECT 42.745 49.965 43.955 51.635 ;
        RECT 42.745 49.425 43.265 52.175 ;
        RECT 40.905 49.945 42.575 51.655 ;
        RECT 40.905 49.425 41.655 52.175 ;
        RECT 35.385 49.945 40.73 51.655 ;
        RECT 35.385 49.425 37.965 52.175 ;
        RECT 29.865 49.945 35.21 51.655 ;
        RECT 29.865 49.425 32.445 52.175 ;
        RECT 29.405 49.99 29.695 51.61 ;
        RECT 28.025 49.965 29.235 51.635 ;
        RECT 28.025 49.425 28.545 52.175 ;
        RECT 26.185 49.945 27.855 51.655 ;
        RECT 26.185 49.425 26.935 52.175 ;
        RECT 20.665 49.945 26.01 51.655 ;
        RECT 20.665 49.425 23.245 52.175 ;
        RECT 15.145 49.945 20.49 51.655 ;
        RECT 15.145 49.425 17.725 52.175 ;
        RECT 14.685 49.99 14.975 51.61 ;
        RECT 13.305 49.965 14.515 51.635 ;
        RECT 13.305 49.425 13.825 52.175 ;
        RECT 10.545 49.945 13.135 51.655 ;
        RECT 10.545 49.425 11.755 52.175 ;
        RECT 10 56.155 189.86 56.325 ;
        RECT 189.025 55.43 189.315 57.05 ;
        RECT 186.265 55.385 188.855 57.095 ;
        RECT 186.265 54.865 187.475 57.615 ;
        RECT 182.585 55.385 186.095 57.095 ;
        RECT 182.585 54.865 184.235 57.615 ;
        RECT 177.065 55.385 182.41 57.095 ;
        RECT 177.065 54.865 179.645 57.615 ;
        RECT 176.605 55.43 176.895 57.05 ;
        RECT 175.225 55.405 176.435 57.075 ;
        RECT 175.225 54.865 175.745 57.615 ;
        RECT 173.385 55.385 175.055 57.095 ;
        RECT 173.385 54.865 174.135 57.615 ;
        RECT 167.865 55.385 173.21 57.095 ;
        RECT 167.865 54.865 170.445 57.615 ;
        RECT 162.345 55.385 167.69 57.095 ;
        RECT 162.345 54.865 164.925 57.615 ;
        RECT 161.885 55.43 162.175 57.05 ;
        RECT 160.505 55.405 161.715 57.075 ;
        RECT 160.505 54.865 161.025 57.615 ;
        RECT 158.665 55.385 160.335 57.095 ;
        RECT 158.665 54.865 159.415 57.615 ;
        RECT 153.145 55.385 158.49 57.095 ;
        RECT 153.145 54.865 155.725 57.615 ;
        RECT 147.625 55.385 152.97 57.095 ;
        RECT 147.625 54.865 150.205 57.615 ;
        RECT 147.165 55.43 147.455 57.05 ;
        RECT 145.785 55.405 146.995 57.075 ;
        RECT 145.785 54.865 146.305 57.615 ;
        RECT 143.945 55.385 145.615 57.095 ;
        RECT 143.945 54.865 144.695 57.615 ;
        RECT 138.425 55.385 143.77 57.095 ;
        RECT 138.425 54.865 141.005 57.615 ;
        RECT 132.905 55.385 138.25 57.095 ;
        RECT 132.905 54.865 135.485 57.615 ;
        RECT 132.445 55.43 132.735 57.05 ;
        RECT 131.065 55.405 132.275 57.075 ;
        RECT 131.065 54.865 131.585 57.615 ;
        RECT 129.225 55.385 130.895 57.095 ;
        RECT 129.225 54.865 129.975 57.615 ;
        RECT 123.705 55.385 129.05 57.095 ;
        RECT 123.705 54.865 126.285 57.615 ;
        RECT 118.185 55.385 123.53 57.095 ;
        RECT 118.185 54.865 120.765 57.615 ;
        RECT 117.725 55.43 118.015 57.05 ;
        RECT 116.345 55.405 117.555 57.075 ;
        RECT 116.345 54.865 116.865 57.615 ;
        RECT 114.505 55.385 116.175 57.095 ;
        RECT 114.505 54.865 115.255 57.615 ;
        RECT 108.985 55.385 114.33 57.095 ;
        RECT 108.985 54.865 111.565 57.615 ;
        RECT 103.465 55.385 108.81 57.095 ;
        RECT 103.465 54.865 106.045 57.615 ;
        RECT 103.005 55.43 103.295 57.05 ;
        RECT 101.625 55.405 102.835 57.075 ;
        RECT 101.625 54.865 102.145 57.615 ;
        RECT 99.785 55.385 101.455 57.095 ;
        RECT 99.785 54.865 100.535 57.615 ;
        RECT 94.265 55.385 99.61 57.095 ;
        RECT 94.265 54.865 96.845 57.615 ;
        RECT 88.745 55.385 94.09 57.095 ;
        RECT 88.745 54.865 91.325 57.615 ;
        RECT 88.285 55.43 88.575 57.05 ;
        RECT 86.905 55.405 88.115 57.075 ;
        RECT 86.905 54.865 87.425 57.615 ;
        RECT 85.065 55.385 86.735 57.095 ;
        RECT 85.065 54.865 85.815 57.615 ;
        RECT 79.545 55.385 84.89 57.095 ;
        RECT 79.545 54.865 82.125 57.615 ;
        RECT 74.025 55.385 79.37 57.095 ;
        RECT 74.025 54.865 76.605 57.615 ;
        RECT 73.565 55.43 73.855 57.05 ;
        RECT 72.185 55.405 73.395 57.075 ;
        RECT 72.185 54.865 72.705 57.615 ;
        RECT 70.345 55.385 72.015 57.095 ;
        RECT 70.345 54.865 71.095 57.615 ;
        RECT 64.825 55.385 70.17 57.095 ;
        RECT 64.825 54.865 67.405 57.615 ;
        RECT 59.305 55.385 64.65 57.095 ;
        RECT 59.305 54.865 61.885 57.615 ;
        RECT 58.845 55.43 59.135 57.05 ;
        RECT 57.465 55.405 58.675 57.075 ;
        RECT 57.465 54.865 57.985 57.615 ;
        RECT 55.625 55.385 57.295 57.095 ;
        RECT 55.625 54.865 56.375 57.615 ;
        RECT 50.105 55.385 55.45 57.095 ;
        RECT 50.105 54.865 52.685 57.615 ;
        RECT 44.585 55.385 49.93 57.095 ;
        RECT 44.585 54.865 47.165 57.615 ;
        RECT 44.125 55.43 44.415 57.05 ;
        RECT 42.745 55.405 43.955 57.075 ;
        RECT 42.745 54.865 43.265 57.615 ;
        RECT 40.905 55.385 42.575 57.095 ;
        RECT 40.905 54.865 41.655 57.615 ;
        RECT 35.385 55.385 40.73 57.095 ;
        RECT 35.385 54.865 37.965 57.615 ;
        RECT 29.865 55.385 35.21 57.095 ;
        RECT 29.865 54.865 32.445 57.615 ;
        RECT 29.405 55.43 29.695 57.05 ;
        RECT 28.025 55.405 29.235 57.075 ;
        RECT 28.025 54.865 28.545 57.615 ;
        RECT 26.185 55.385 27.855 57.095 ;
        RECT 26.185 54.865 26.935 57.615 ;
        RECT 20.665 55.385 26.01 57.095 ;
        RECT 20.665 54.865 23.245 57.615 ;
        RECT 15.145 55.385 20.49 57.095 ;
        RECT 15.145 54.865 17.725 57.615 ;
        RECT 14.685 55.43 14.975 57.05 ;
        RECT 13.305 55.405 14.515 57.075 ;
        RECT 13.305 54.865 13.825 57.615 ;
        RECT 10.545 55.385 13.135 57.095 ;
        RECT 10.545 54.865 11.755 57.615 ;
        RECT 10 12.635 189.86 12.805 ;
        RECT 189.025 11.91 189.315 13.53 ;
        RECT 186.265 11.865 188.855 13.575 ;
        RECT 186.265 11.345 187.475 14.095 ;
        RECT 182.585 11.865 186.095 13.575 ;
        RECT 182.585 11.345 184.235 14.095 ;
        RECT 177.065 11.865 182.41 13.575 ;
        RECT 177.065 11.345 179.645 14.095 ;
        RECT 176.605 11.91 176.895 13.53 ;
        RECT 175.225 11.885 176.435 13.555 ;
        RECT 175.225 11.345 175.745 14.095 ;
        RECT 172.465 11.865 175.055 13.575 ;
        RECT 172.465 11.345 173.675 13.575 ;
        RECT 171.545 12.635 173.195 14.095 ;
        RECT 168.785 11.865 172.295 12.805 ;
        RECT 170.615 11.865 170.945 13.285 ;
        RECT 168.785 11.345 170.435 12.805 ;
        RECT 168.355 12.635 168.685 13.285 ;
        RECT 167.895 11.835 168.225 12.805 ;
        RECT 162.345 12.635 167.69 13.575 ;
        RECT 167.055 12.155 167.385 13.575 ;
        RECT 166.215 12.155 166.545 13.575 ;
        RECT 165.375 12.155 165.705 13.575 ;
        RECT 162.345 12.635 164.925 14.095 ;
        RECT 164.535 12.155 164.865 14.095 ;
        RECT 163.695 12.155 164.025 14.095 ;
        RECT 161.885 11.91 162.175 13.53 ;
        RECT 160.505 11.885 161.715 13.555 ;
        RECT 160.505 11.345 161.025 14.095 ;
        RECT 158.665 11.865 160.335 13.575 ;
        RECT 158.665 11.865 159.415 14.095 ;
        RECT 157.745 11.345 158.955 12.805 ;
        RECT 153.145 12.635 158.49 13.575 ;
        RECT 154.065 11.865 157.575 13.575 ;
        RECT 153.145 12.635 155.725 14.095 ;
        RECT 154.065 11.345 155.715 14.095 ;
        RECT 153.175 11.835 153.505 14.095 ;
        RECT 147.625 12.635 152.97 13.575 ;
        RECT 152.335 12.155 152.665 13.575 ;
        RECT 151.495 12.155 151.825 13.575 ;
        RECT 150.655 12.155 150.985 13.575 ;
        RECT 147.625 12.635 150.205 14.095 ;
        RECT 149.815 12.155 150.145 14.095 ;
        RECT 148.975 12.155 149.305 14.095 ;
        RECT 147.165 11.91 147.455 13.53 ;
        RECT 145.785 11.885 146.995 12.805 ;
        RECT 145.785 11.345 146.305 12.805 ;
        RECT 144.865 12.635 146.075 13.555 ;
        RECT 143.945 11.865 145.615 12.805 ;
        RECT 144.865 11.865 145.385 14.095 ;
        RECT 143.945 11.345 144.695 12.805 ;
        RECT 143.935 12.635 144.265 13.285 ;
        RECT 143.095 12.635 143.425 13.285 ;
        RECT 143.055 11.835 143.385 12.805 ;
        RECT 142.255 12.635 142.585 13.285 ;
        RECT 142.215 12.155 142.545 12.805 ;
        RECT 141.415 12.635 141.745 13.285 ;
        RECT 141.375 12.155 141.705 12.805 ;
        RECT 140.575 12.635 140.905 13.285 ;
        RECT 140.535 12.155 140.865 12.805 ;
        RECT 139.735 12.635 140.065 13.605 ;
        RECT 139.695 12.155 140.025 12.805 ;
        RECT 138.855 12.155 139.185 12.805 ;
        RECT 132.905 11.865 138.25 12.805 ;
        RECT 137.535 11.865 137.865 13.605 ;
        RECT 136.695 11.865 137.025 13.285 ;
        RECT 135.855 11.865 136.185 13.285 ;
        RECT 132.905 11.345 135.485 12.805 ;
        RECT 135.015 11.345 135.345 13.285 ;
        RECT 134.175 11.345 134.505 13.285 ;
        RECT 133.335 11.345 133.665 13.285 ;
        RECT 132.445 11.91 132.735 13.53 ;
        RECT 131.065 11.885 132.275 13.555 ;
        RECT 131.065 11.345 131.585 14.095 ;
        RECT 127.385 12.635 130.895 13.575 ;
        RECT 129.225 11.865 130.895 13.575 ;
        RECT 129.225 11.345 129.975 13.575 ;
        RECT 123.705 11.865 129.05 12.805 ;
        RECT 127.385 11.865 129.035 14.095 ;
        RECT 121.865 12.635 127.21 13.575 ;
        RECT 123.705 11.345 126.285 13.575 ;
        RECT 121.865 12.635 124.445 14.095 ;
        RECT 122.775 12.155 123.105 14.095 ;
        RECT 121.935 12.155 122.265 14.095 ;
        RECT 121.095 12.155 121.425 12.805 ;
        RECT 120.875 12.635 121.205 13.285 ;
        RECT 120.255 12.155 120.585 12.805 ;
        RECT 119.415 12.155 119.745 12.805 ;
        RECT 118.615 12.635 118.945 13.285 ;
        RECT 118.575 11.835 118.905 12.805 ;
        RECT 117.725 11.91 118.015 13.53 ;
        RECT 116.345 11.885 117.555 13.575 ;
        RECT 116.345 11.345 116.865 13.575 ;
        RECT 115.885 12.635 116.635 14.095 ;
        RECT 114.505 11.865 116.175 12.805 ;
        RECT 114.955 11.865 115.285 13.285 ;
        RECT 114.505 11.345 115.255 12.805 ;
        RECT 114.115 12.635 114.445 13.285 ;
        RECT 108.985 11.865 114.33 12.805 ;
        RECT 113.275 11.865 113.605 13.285 ;
        RECT 112.435 11.865 112.765 13.285 ;
        RECT 111.595 11.865 111.925 13.285 ;
        RECT 108.985 11.345 111.565 12.805 ;
        RECT 110.755 11.345 111.085 13.605 ;
        RECT 108.985 11.345 110.195 13.555 ;
        RECT 108.985 11.345 109.505 14.095 ;
        RECT 103.465 11.865 108.81 12.805 ;
        RECT 108.095 11.865 108.425 13.605 ;
        RECT 107.255 11.865 107.585 13.285 ;
        RECT 106.415 11.865 106.745 13.285 ;
        RECT 103.465 11.345 106.045 12.805 ;
        RECT 105.575 11.345 105.905 13.285 ;
        RECT 104.735 11.345 105.065 13.285 ;
        RECT 103.895 11.345 104.225 13.285 ;
        RECT 103.005 11.91 103.295 13.53 ;
        RECT 100.245 12.635 102.835 13.575 ;
        RECT 102.115 11.835 102.445 13.575 ;
        RECT 101.275 12.155 101.605 13.575 ;
        RECT 100.245 12.635 101.455 14.095 ;
        RECT 100.435 12.155 100.765 14.095 ;
        RECT 96.565 12.635 100.075 13.575 ;
        RECT 99.595 12.155 99.925 13.575 ;
        RECT 98.755 12.155 99.085 13.575 ;
        RECT 97.915 12.155 98.245 13.575 ;
        RECT 96.565 12.635 98.215 14.095 ;
        RECT 96.135 11.835 96.465 12.805 ;
        RECT 95.575 12.635 95.905 13.285 ;
        RECT 95.295 12.155 95.625 12.805 ;
        RECT 94.455 12.155 94.785 12.805 ;
        RECT 93.615 12.155 93.945 12.805 ;
        RECT 93.315 12.635 93.645 13.285 ;
        RECT 92.775 12.155 93.105 12.805 ;
        RECT 91.505 12.635 92.715 13.555 ;
        RECT 91.935 12.155 92.265 13.555 ;
        RECT 91.505 12.635 92.025 14.095 ;
        RECT 88.745 11.865 91.335 13.575 ;
        RECT 88.745 11.345 89.955 14.095 ;
        RECT 88.285 11.91 88.575 13.53 ;
        RECT 86.905 12.635 88.115 13.555 ;
        RECT 87.395 11.835 87.725 13.555 ;
        RECT 86.905 12.635 87.425 14.095 ;
        RECT 86.555 12.155 86.885 12.805 ;
        RECT 85.065 12.635 86.735 13.575 ;
        RECT 85.715 12.155 86.045 13.575 ;
        RECT 85.065 12.635 85.815 14.095 ;
        RECT 84.875 12.155 85.205 12.805 ;
        RECT 79.545 12.635 84.89 13.575 ;
        RECT 84.035 12.155 84.365 13.575 ;
        RECT 83.195 12.155 83.525 13.575 ;
        RECT 81.385 11.885 82.595 13.575 ;
        RECT 79.545 12.635 82.125 14.095 ;
        RECT 81.385 11.345 81.905 14.095 ;
        RECT 79.545 11.865 81.215 14.095 ;
        RECT 79.545 11.345 80.295 14.095 ;
        RECT 74.025 12.635 79.37 13.575 ;
        RECT 78.655 11.835 78.985 13.575 ;
        RECT 77.815 12.155 78.145 13.575 ;
        RECT 76.975 12.155 77.305 13.575 ;
        RECT 74.025 12.635 76.605 14.095 ;
        RECT 76.135 12.155 76.465 14.095 ;
        RECT 75.295 12.155 75.625 14.095 ;
        RECT 74.455 12.155 74.785 14.095 ;
        RECT 73.565 11.91 73.855 13.53 ;
        RECT 68.045 11.865 73.39 12.805 ;
        RECT 71.265 11.865 72.475 13.555 ;
        RECT 71.265 11.865 71.785 14.095 ;
        RECT 70.375 11.865 70.705 13.605 ;
        RECT 68.045 11.345 70.625 12.805 ;
        RECT 69.535 11.345 69.865 13.285 ;
        RECT 68.695 11.345 69.025 13.285 ;
        RECT 67.855 12.635 68.185 13.285 ;
        RECT 67.155 11.835 67.485 12.805 ;
        RECT 67.015 12.635 67.345 13.285 ;
        RECT 66.315 12.155 66.645 12.805 ;
        RECT 66.175 12.635 66.505 13.285 ;
        RECT 65.475 12.155 65.805 12.805 ;
        RECT 64.365 12.635 65.575 13.555 ;
        RECT 64.635 12.155 64.965 13.555 ;
        RECT 64.365 12.635 64.885 14.095 ;
        RECT 63.795 12.155 64.125 12.805 ;
        RECT 63.435 12.635 63.765 13.285 ;
        RECT 62.955 12.155 63.285 12.805 ;
        RECT 61.145 11.885 62.355 12.805 ;
        RECT 61.145 11.345 61.665 12.805 ;
        RECT 61.175 11.345 61.505 13.285 ;
        RECT 59.305 11.865 60.975 12.805 ;
        RECT 59.305 11.865 60.515 13.555 ;
        RECT 59.305 11.345 60.055 13.555 ;
        RECT 59.305 11.345 59.825 14.095 ;
        RECT 58.845 11.91 59.135 13.53 ;
        RECT 57.005 12.635 58.675 13.575 ;
        RECT 53.325 11.865 58.67 12.805 ;
        RECT 57.005 11.865 57.755 14.095 ;
        RECT 54.245 11.865 56.835 13.575 ;
        RECT 53.325 11.345 55.905 12.805 ;
        RECT 54.245 11.345 55.455 14.095 ;
        RECT 53.255 12.635 53.585 13.285 ;
        RECT 52.435 11.835 52.765 12.805 ;
        RECT 51.595 12.155 51.925 12.805 ;
        RECT 50.995 12.635 51.325 13.285 ;
        RECT 50.755 12.155 51.085 12.805 ;
        RECT 47.805 12.635 50.395 13.575 ;
        RECT 49.915 12.155 50.245 13.575 ;
        RECT 49.075 12.155 49.405 13.575 ;
        RECT 47.805 12.635 49.015 14.095 ;
        RECT 48.235 12.155 48.565 14.095 ;
        RECT 46.425 11.885 47.635 12.805 ;
        RECT 46.785 11.885 47.165 13.205 ;
        RECT 46.425 11.345 46.945 12.805 ;
        RECT 45.945 12.635 46.275 13.205 ;
        RECT 44.585 11.865 46.255 12.805 ;
        RECT 44.585 11.345 45.335 12.805 ;
        RECT 44.125 11.91 44.415 13.53 ;
        RECT 42.745 11.885 43.955 13.555 ;
        RECT 42.745 11.345 43.265 14.095 ;
        RECT 40.905 11.865 42.575 13.575 ;
        RECT 40.905 11.345 41.655 14.095 ;
        RECT 38.145 12.635 40.735 13.575 ;
        RECT 35.385 11.865 40.73 12.805 ;
        RECT 38.145 11.865 39.355 14.095 ;
        RECT 35.385 11.345 37.965 12.805 ;
        RECT 37.215 11.345 37.545 13.285 ;
        RECT 36.375 11.345 36.705 13.285 ;
        RECT 35.535 11.345 35.865 13.285 ;
        RECT 34.695 12.635 35.025 13.285 ;
        RECT 34.495 11.835 34.825 12.805 ;
        RECT 33.855 12.635 34.185 13.285 ;
        RECT 33.655 12.155 33.985 12.805 ;
        RECT 33.015 12.635 33.345 13.605 ;
        RECT 32.815 12.155 33.145 12.805 ;
        RECT 29.865 12.635 32.455 13.575 ;
        RECT 31.975 12.155 32.305 13.575 ;
        RECT 31.135 12.155 31.465 13.575 ;
        RECT 29.865 12.635 31.075 14.095 ;
        RECT 30.295 12.155 30.625 14.095 ;
        RECT 29.405 11.91 29.695 13.53 ;
        RECT 28.025 11.885 29.235 13.575 ;
        RECT 28.025 11.345 28.545 13.575 ;
        RECT 27.565 12.635 28.315 14.095 ;
        RECT 26.185 11.865 27.855 12.805 ;
        RECT 24.805 12.635 27.395 13.575 ;
        RECT 26.185 11.345 26.935 13.575 ;
        RECT 24.805 12.635 26.015 14.095 ;
        RECT 20.665 11.865 26.01 12.805 ;
        RECT 23.915 11.865 24.245 13.605 ;
        RECT 23.075 11.865 23.405 13.285 ;
        RECT 20.665 11.345 23.245 12.805 ;
        RECT 22.235 11.345 22.565 13.285 ;
        RECT 21.395 11.345 21.725 13.285 ;
        RECT 20.555 12.635 20.885 13.285 ;
        RECT 15.145 11.865 20.49 12.805 ;
        RECT 19.715 11.865 20.045 13.285 ;
        RECT 17.905 11.865 19.115 13.555 ;
        RECT 17.905 11.865 18.425 14.095 ;
        RECT 15.145 11.865 17.735 13.575 ;
        RECT 15.145 11.345 17.725 13.575 ;
        RECT 15.145 11.345 16.355 14.095 ;
        RECT 14.685 11.91 14.975 13.53 ;
        RECT 13.305 11.885 14.515 13.555 ;
        RECT 13.305 11.345 13.825 14.095 ;
        RECT 10.545 11.865 13.135 13.575 ;
        RECT 10.545 11.345 11.755 14.095 ;
        RECT 10 18.075 189.86 18.245 ;
        RECT 189.025 17.35 189.315 18.97 ;
        RECT 186.265 17.305 188.855 19.015 ;
        RECT 186.265 16.785 187.475 19.535 ;
        RECT 182.585 17.305 186.095 19.015 ;
        RECT 182.585 16.785 184.235 19.535 ;
        RECT 177.065 18.075 182.41 19.015 ;
        RECT 181.695 17.275 182.025 19.015 ;
        RECT 180.855 17.595 181.185 19.015 ;
        RECT 180.015 17.595 180.345 19.015 ;
        RECT 177.065 18.075 179.645 19.535 ;
        RECT 179.175 17.595 179.505 19.535 ;
        RECT 178.335 17.595 178.665 19.535 ;
        RECT 177.495 17.595 177.825 19.535 ;
        RECT 176.605 17.35 176.895 18.97 ;
        RECT 174.765 18.075 176.435 19.015 ;
        RECT 175.715 17.465 175.885 19.015 ;
        RECT 174.765 18.075 175.515 19.535 ;
        RECT 174.745 17.545 174.955 18.245 ;
        RECT 174.255 18.075 174.59 18.645 ;
        RECT 173.395 18.075 173.67 18.725 ;
        RECT 172.56 17.575 172.93 18.245 ;
        RECT 172.035 18.075 172.205 18.855 ;
        RECT 171.065 18.075 171.275 18.775 ;
        RECT 170.615 17.615 170.865 18.245 ;
        RECT 169.675 17.695 170.005 18.245 ;
        RECT 168.88 18.075 169.25 18.745 ;
        RECT 167.865 17.325 169.075 18.245 ;
        RECT 167.865 16.785 168.385 18.245 ;
        RECT 166.975 17.275 167.305 18.245 ;
        RECT 166.935 18.075 167.185 18.705 ;
        RECT 166.135 17.595 166.465 18.245 ;
        RECT 165.995 18.075 166.325 18.625 ;
        RECT 165.295 17.595 165.625 18.245 ;
        RECT 164.455 17.595 164.785 18.245 ;
        RECT 164.335 18.075 164.66 18.705 ;
        RECT 163.615 17.595 163.945 18.245 ;
        RECT 162.915 18.075 163.185 18.705 ;
        RECT 162.775 17.595 163.105 18.245 ;
        RECT 161.885 17.35 162.175 18.97 ;
        RECT 160.505 18.075 161.715 18.995 ;
        RECT 160.505 18.075 161.025 19.535 ;
        RECT 160.075 17.465 160.245 18.245 ;
        RECT 159.615 18.075 159.785 18.855 ;
        RECT 159.105 17.545 159.315 18.245 ;
        RECT 158.645 18.075 158.855 18.775 ;
        RECT 156.92 17.575 157.29 18.245 ;
        RECT 156.46 18.075 156.83 18.745 ;
        RECT 154.975 17.615 155.225 18.245 ;
        RECT 154.515 18.075 154.765 18.705 ;
        RECT 154.035 17.695 154.365 18.245 ;
        RECT 153.575 18.075 153.905 18.625 ;
        RECT 152.225 17.325 153.435 18.245 ;
        RECT 147.625 18.075 152.97 19.015 ;
        RECT 152.225 16.785 152.745 19.015 ;
        RECT 150.385 17.305 152.055 19.015 ;
        RECT 150.385 16.785 151.135 19.015 ;
        RECT 147.625 17.305 150.215 19.015 ;
        RECT 147.625 17.305 150.205 19.535 ;
        RECT 147.625 16.785 148.835 19.535 ;
        RECT 147.165 17.35 147.455 18.97 ;
        RECT 145.255 17.595 145.585 18.725 ;
        RECT 142.995 17.595 143.325 18.725 ;
        RECT 141.185 17.325 142.395 18.245 ;
        RECT 141.185 16.785 141.705 18.245 ;
        RECT 140.265 18.075 141.475 18.995 ;
        RECT 138.425 17.305 141.015 18.245 ;
        RECT 140.265 17.305 140.785 19.535 ;
        RECT 138.425 16.785 139.635 18.245 ;
        RECT 139.375 16.785 139.545 18.855 ;
        RECT 138.405 18.075 138.615 18.775 ;
        RECT 137.435 17.595 137.765 18.245 ;
        RECT 136.22 18.075 136.59 18.745 ;
        RECT 135.175 17.595 135.505 18.245 ;
        RECT 132.905 17.305 134.575 18.245 ;
        RECT 134.275 17.305 134.525 18.705 ;
        RECT 133.335 17.305 133.665 18.625 ;
        RECT 132.905 16.785 133.655 18.245 ;
        RECT 132.445 17.35 132.735 18.97 ;
        RECT 131.065 17.325 132.275 18.995 ;
        RECT 131.065 16.785 131.585 19.535 ;
        RECT 129.225 17.305 130.895 18.245 ;
        RECT 125.545 18.075 130.89 19.015 ;
        RECT 129.225 16.785 129.975 19.015 ;
        RECT 128.235 17.595 128.565 19.015 ;
        RECT 125.545 18.075 128.125 19.535 ;
        RECT 125.975 17.595 126.305 19.535 ;
        RECT 123.705 17.305 125.375 18.245 ;
        RECT 124.655 17.305 124.825 18.855 ;
        RECT 123.705 16.785 124.455 18.245 ;
        RECT 123.685 18.075 123.895 18.775 ;
        RECT 122.775 17.595 123.105 18.245 ;
        RECT 121.935 17.595 122.265 18.245 ;
        RECT 121.5 18.075 121.87 18.745 ;
        RECT 121.095 17.595 121.425 18.245 ;
        RECT 120.255 17.595 120.585 18.245 ;
        RECT 119.555 18.075 119.805 18.705 ;
        RECT 119.415 17.595 119.745 18.245 ;
        RECT 118.615 18.075 118.945 18.625 ;
        RECT 118.575 17.275 118.905 18.245 ;
        RECT 117.725 17.35 118.015 18.97 ;
        RECT 114.965 17.305 117.555 19.015 ;
        RECT 114.965 16.785 116.175 19.535 ;
        RECT 114.035 18.075 114.365 18.725 ;
        RECT 113.975 17.595 114.305 18.245 ;
        RECT 113.195 18.075 113.525 18.725 ;
        RECT 112.355 18.075 112.685 18.725 ;
        RECT 111.715 17.595 112.045 18.245 ;
        RECT 111.515 18.075 111.845 18.725 ;
        RECT 110.675 18.075 111.005 18.725 ;
        RECT 108.985 17.325 110.195 18.245 ;
        RECT 109.835 17.325 110.165 19.045 ;
        RECT 108.985 16.785 109.505 18.245 ;
        RECT 108.065 18.075 109.275 18.995 ;
        RECT 108.065 18.075 108.585 19.535 ;
        RECT 108.095 17.275 108.425 19.535 ;
        RECT 106.225 18.075 107.895 19.015 ;
        RECT 107.255 17.595 107.585 19.015 ;
        RECT 106.225 18.075 106.975 19.535 ;
        RECT 106.415 17.595 106.745 19.535 ;
        RECT 103.465 18.075 106.055 19.015 ;
        RECT 105.575 17.595 105.905 19.015 ;
        RECT 104.735 17.595 105.065 19.015 ;
        RECT 103.465 18.075 104.675 19.535 ;
        RECT 103.895 17.595 104.225 19.535 ;
        RECT 103.005 17.35 103.295 18.97 ;
        RECT 101.165 17.305 102.835 19.015 ;
        RECT 101.165 16.785 101.915 19.535 ;
        RECT 98.405 17.305 100.995 18.245 ;
        RECT 100.275 17.305 100.445 18.855 ;
        RECT 98.405 16.785 99.615 18.245 ;
        RECT 99.305 16.785 99.515 18.775 ;
        RECT 97.475 17.595 97.805 18.245 ;
        RECT 97.12 18.075 97.49 18.745 ;
        RECT 95.215 17.595 95.545 18.245 ;
        RECT 95.175 18.075 95.425 18.705 ;
        RECT 94.235 18.075 94.565 18.625 ;
        RECT 93.345 17.325 94.555 18.245 ;
        RECT 93.345 16.785 93.865 18.245 ;
        RECT 92.425 18.075 93.635 18.995 ;
        RECT 91.505 17.305 93.175 18.245 ;
        RECT 92.425 17.305 92.945 19.535 ;
        RECT 88.745 18.075 92.255 19.015 ;
        RECT 91.505 16.785 92.255 19.015 ;
        RECT 88.745 17.305 91.335 19.015 ;
        RECT 88.745 17.305 90.395 19.535 ;
        RECT 88.745 16.785 89.955 19.535 ;
        RECT 88.285 17.35 88.575 18.97 ;
        RECT 86.905 17.325 88.115 19.015 ;
        RECT 86.905 16.785 87.425 19.015 ;
        RECT 86.445 18.075 87.195 19.535 ;
        RECT 85.065 17.305 86.735 18.245 ;
        RECT 85.065 16.785 85.815 18.245 ;
        RECT 85.455 16.785 85.785 18.725 ;
        RECT 84.135 17.595 84.465 18.245 ;
        RECT 83.195 18.075 83.525 18.725 ;
        RECT 81.875 17.595 82.205 18.245 ;
        RECT 81.875 17.595 82.045 18.855 ;
        RECT 79.545 17.305 81.215 18.245 ;
        RECT 80.905 17.305 81.115 18.775 ;
        RECT 79.545 16.785 80.295 18.245 ;
        RECT 78.72 18.075 79.09 18.745 ;
        RECT 78.655 17.275 78.985 18.245 ;
        RECT 77.815 17.595 78.145 18.245 ;
        RECT 76.975 17.595 77.305 18.245 ;
        RECT 76.775 18.075 77.025 18.705 ;
        RECT 76.135 17.595 76.465 18.245 ;
        RECT 75.835 18.075 76.165 18.625 ;
        RECT 75.295 17.595 75.625 18.245 ;
        RECT 74.025 18.075 75.235 18.995 ;
        RECT 74.455 17.595 74.785 18.995 ;
        RECT 74.025 18.075 74.545 19.535 ;
        RECT 73.565 17.35 73.855 18.97 ;
        RECT 72.185 17.325 73.395 18.995 ;
        RECT 72.185 16.785 72.705 19.535 ;
        RECT 71.255 17.595 71.585 18.725 ;
        RECT 68.995 17.595 69.325 18.725 ;
        RECT 66.665 17.305 68.335 19.015 ;
        RECT 66.665 16.785 67.415 19.535 ;
        RECT 65.775 17.465 65.945 18.855 ;
        RECT 64.805 17.545 65.015 18.775 ;
        RECT 62.62 17.575 62.99 18.745 ;
        RECT 60.675 17.615 60.925 18.705 ;
        RECT 59.735 17.695 60.065 18.625 ;
        RECT 58.845 17.35 59.135 18.97 ;
        RECT 57.465 17.325 58.675 19.015 ;
        RECT 57.465 16.785 57.985 19.015 ;
        RECT 57.005 18.075 57.755 19.535 ;
        RECT 56.575 17.465 56.745 18.245 ;
        RECT 56.115 18.075 56.285 18.855 ;
        RECT 55.605 17.545 55.815 18.245 ;
        RECT 55.145 18.075 55.355 18.775 ;
        RECT 53.42 17.575 53.79 18.245 ;
        RECT 52.96 18.075 53.33 18.745 ;
        RECT 51.475 17.615 51.725 18.245 ;
        RECT 51.015 18.075 51.265 18.705 ;
        RECT 50.535 17.695 50.865 18.245 ;
        RECT 50.075 18.075 50.405 18.625 ;
        RECT 48.265 17.305 49.935 18.245 ;
        RECT 48.265 17.305 49.475 18.995 ;
        RECT 48.265 16.785 49.015 18.995 ;
        RECT 48.265 16.785 48.785 19.535 ;
        RECT 44.585 18.075 48.095 19.015 ;
        RECT 47.275 17.595 47.605 19.015 ;
        RECT 44.585 18.075 46.235 19.535 ;
        RECT 45.015 17.595 45.345 19.535 ;
        RECT 44.125 17.35 44.415 18.97 ;
        RECT 42.745 17.305 43.955 18.995 ;
        RECT 42.745 17.305 43.265 19.535 ;
        RECT 41.365 17.305 43.955 18.245 ;
        RECT 41.365 16.785 42.575 19.015 ;
        RECT 40.905 18.075 41.655 19.535 ;
        RECT 40.435 17.595 40.765 18.245 ;
        RECT 35.385 18.075 40.73 19.015 ;
        RECT 39.595 17.595 39.925 19.015 ;
        RECT 38.755 17.595 39.085 19.015 ;
        RECT 37.915 17.595 38.245 19.015 ;
        RECT 35.385 18.075 37.965 19.535 ;
        RECT 37.075 17.595 37.405 19.535 ;
        RECT 36.235 17.275 36.565 19.535 ;
        RECT 29.865 18.075 35.21 19.015 ;
        RECT 34.495 17.275 34.825 19.015 ;
        RECT 33.655 17.595 33.985 19.015 ;
        RECT 32.815 17.595 33.145 19.015 ;
        RECT 29.865 18.075 32.445 19.535 ;
        RECT 31.975 17.595 32.305 19.535 ;
        RECT 31.135 17.595 31.465 19.535 ;
        RECT 30.295 17.595 30.625 19.535 ;
        RECT 29.405 17.35 29.695 18.97 ;
        RECT 28.025 17.305 29.235 18.995 ;
        RECT 28.025 17.305 28.545 19.535 ;
        RECT 27.565 16.785 28.315 18.245 ;
        RECT 26.185 18.075 27.855 19.015 ;
        RECT 24.805 17.305 27.395 18.245 ;
        RECT 26.185 17.305 26.935 19.535 ;
        RECT 24.805 16.785 26.015 18.245 ;
        RECT 20.665 18.075 26.01 19.015 ;
        RECT 23.915 17.275 24.245 19.015 ;
        RECT 23.075 17.595 23.405 19.015 ;
        RECT 20.665 18.075 23.245 19.535 ;
        RECT 22.235 17.595 22.565 19.535 ;
        RECT 21.395 17.595 21.725 19.535 ;
        RECT 20.555 17.595 20.885 18.245 ;
        RECT 15.145 18.075 20.49 19.015 ;
        RECT 19.715 17.595 20.045 19.015 ;
        RECT 17.905 17.325 19.115 19.015 ;
        RECT 17.905 16.785 18.425 19.015 ;
        RECT 15.145 17.305 17.735 19.015 ;
        RECT 15.145 17.305 17.725 19.535 ;
        RECT 15.145 16.785 16.355 19.535 ;
        RECT 14.685 17.35 14.975 18.97 ;
        RECT 13.305 17.325 14.515 18.995 ;
        RECT 13.305 16.785 13.825 19.535 ;
        RECT 10.545 17.305 13.135 19.015 ;
        RECT 10.545 16.785 11.755 19.535 ;
        RECT 10 23.515 189.86 23.685 ;
        RECT 189.025 22.79 189.315 24.41 ;
        RECT 187.645 22.745 188.855 24.435 ;
        RECT 187.645 22.745 188.165 24.975 ;
        RECT 187.185 22.225 187.935 23.685 ;
        RECT 185.805 23.515 187.475 24.455 ;
        RECT 184.425 22.745 187.015 23.685 ;
        RECT 185.805 22.745 186.555 24.975 ;
        RECT 184.425 22.225 185.635 23.685 ;
        RECT 184.915 22.225 185.245 24.485 ;
        RECT 184.075 23.515 184.405 24.165 ;
        RECT 183.535 22.905 183.705 23.685 ;
        RECT 183.235 23.515 183.565 24.165 ;
        RECT 182.565 22.985 182.775 23.685 ;
        RECT 182.395 23.515 182.725 24.165 ;
        RECT 181.555 23.515 181.885 24.165 ;
        RECT 180.715 23.515 181.045 24.165 ;
        RECT 180.38 23.015 180.75 23.685 ;
        RECT 178.905 23.515 180.115 24.435 ;
        RECT 178.905 23.515 179.425 24.975 ;
        RECT 177.065 23.515 178.735 24.455 ;
        RECT 178.435 23.055 178.685 24.455 ;
        RECT 177.495 23.135 177.825 24.455 ;
        RECT 177.065 23.515 177.815 24.975 ;
        RECT 176.605 22.79 176.895 24.41 ;
        RECT 175.225 22.765 176.435 24.455 ;
        RECT 175.225 22.225 175.745 24.455 ;
        RECT 174.765 23.515 175.515 24.975 ;
        RECT 173.385 22.745 175.055 23.685 ;
        RECT 172.005 23.515 174.595 24.455 ;
        RECT 173.385 22.225 174.135 24.455 ;
        RECT 172.005 23.515 173.215 24.975 ;
        RECT 172.875 23.115 173.21 24.975 ;
        RECT 172.015 23.035 172.29 24.975 ;
        RECT 171.525 23.515 171.815 24.415 ;
        RECT 170.605 23.135 170.935 23.685 ;
        RECT 169.775 23.515 170.445 24.055 ;
        RECT 167.865 23.515 169.075 24.435 ;
        RECT 168.815 22.905 168.985 24.435 ;
        RECT 167.865 23.515 168.385 24.975 ;
        RECT 167.845 22.985 168.055 23.685 ;
        RECT 162.345 23.515 167.69 24.455 ;
        RECT 165.66 23.015 166.03 24.455 ;
        RECT 162.345 23.515 164.925 24.975 ;
        RECT 163.715 23.055 163.965 24.975 ;
        RECT 162.775 23.135 163.105 24.975 ;
        RECT 161.885 22.79 162.175 24.41 ;
        RECT 160.505 23.515 161.715 24.435 ;
        RECT 160.505 23.515 161.025 24.975 ;
        RECT 158.665 23.515 160.335 24.455 ;
        RECT 160.075 22.905 160.245 24.455 ;
        RECT 158.665 23.515 159.415 24.975 ;
        RECT 159.105 22.985 159.315 24.975 ;
        RECT 157.735 23.515 158.065 24.165 ;
        RECT 156.92 23.015 157.29 23.685 ;
        RECT 155.475 23.515 155.805 24.165 ;
        RECT 154.975 23.055 155.225 23.685 ;
        RECT 153.145 23.515 154.815 24.455 ;
        RECT 154.035 23.135 154.365 24.455 ;
        RECT 153.145 23.515 153.895 24.975 ;
        RECT 152.225 22.765 153.435 23.685 ;
        RECT 152.225 22.225 152.745 23.685 ;
        RECT 152.215 23.515 152.545 24.165 ;
        RECT 150.385 22.745 152.055 23.685 ;
        RECT 151.375 22.745 151.705 24.165 ;
        RECT 150.385 22.225 151.135 23.685 ;
        RECT 150.535 22.225 150.865 24.165 ;
        RECT 147.625 22.745 150.215 23.685 ;
        RECT 149.695 22.745 150.025 24.165 ;
        RECT 148.855 22.745 149.185 24.165 ;
        RECT 147.625 22.225 148.835 23.685 ;
        RECT 148.015 22.225 148.345 24.485 ;
        RECT 147.165 22.79 147.455 24.41 ;
        RECT 145.785 22.765 146.995 23.685 ;
        RECT 141.645 23.515 146.99 24.455 ;
        RECT 145.785 22.225 146.305 24.455 ;
        RECT 142.105 22.745 145.615 24.455 ;
        RECT 141.645 23.515 144.225 24.975 ;
        RECT 142.105 22.225 143.755 24.975 ;
        RECT 141.215 22.905 141.385 23.685 ;
        RECT 140.715 23.515 141.045 24.165 ;
        RECT 140.245 22.985 140.455 23.685 ;
        RECT 138.455 23.515 138.785 24.165 ;
        RECT 138.06 23.015 138.43 23.685 ;
        RECT 136.585 23.515 137.795 24.435 ;
        RECT 136.585 23.515 137.105 24.975 ;
        RECT 132.905 23.515 136.415 24.455 ;
        RECT 136.115 23.055 136.365 24.455 ;
        RECT 135.175 23.135 135.505 24.455 ;
        RECT 132.905 23.515 134.555 24.975 ;
        RECT 133.805 23.135 134.135 24.975 ;
        RECT 132.445 22.79 132.735 24.41 ;
        RECT 131.065 23.515 132.275 24.435 ;
        RECT 131.065 23.515 131.585 24.975 ;
        RECT 131.095 22.905 131.265 24.975 ;
        RECT 125.545 23.515 130.89 24.455 ;
        RECT 130.125 22.985 130.335 24.455 ;
        RECT 127.94 23.015 128.31 24.455 ;
        RECT 125.545 23.515 128.125 24.975 ;
        RECT 125.995 23.055 126.245 24.975 ;
        RECT 125.055 23.135 125.385 23.685 ;
        RECT 124.655 23.515 124.825 24.295 ;
        RECT 121.865 22.745 124.455 23.685 ;
        RECT 123.685 22.745 123.895 24.215 ;
        RECT 121.865 22.225 123.075 23.685 ;
        RECT 121.5 23.515 121.87 24.185 ;
        RECT 118.185 22.745 121.695 23.685 ;
        RECT 118.185 22.225 119.835 23.685 ;
        RECT 119.555 22.225 119.805 24.145 ;
        RECT 118.615 22.225 118.945 24.065 ;
        RECT 117.725 22.79 118.015 24.41 ;
        RECT 116.345 23.515 117.555 24.435 ;
        RECT 116.835 22.905 117.005 24.435 ;
        RECT 116.345 23.515 116.865 24.975 ;
        RECT 115.865 22.985 116.075 23.685 ;
        RECT 115.355 23.515 115.685 24.165 ;
        RECT 113.68 23.015 114.05 23.685 ;
        RECT 113.095 23.515 113.425 24.165 ;
        RECT 108.985 23.515 112.495 24.455 ;
        RECT 111.735 23.055 111.985 24.455 ;
        RECT 110.795 23.135 111.125 24.455 ;
        RECT 108.985 23.515 110.635 24.975 ;
        RECT 108.985 22.765 110.195 24.975 ;
        RECT 108.985 22.225 109.505 24.975 ;
        RECT 103.465 22.745 108.81 24.455 ;
        RECT 103.465 22.225 106.045 24.975 ;
        RECT 103.005 22.79 103.295 24.41 ;
        RECT 101.165 23.515 102.835 24.455 ;
        RECT 102.115 22.905 102.285 24.455 ;
        RECT 101.165 23.515 101.915 24.975 ;
        RECT 101.145 22.985 101.355 23.685 ;
        RECT 98.405 23.515 100.995 24.455 ;
        RECT 98.405 23.515 99.615 24.975 ;
        RECT 98.96 23.015 99.33 24.975 ;
        RECT 97.515 23.515 97.685 24.295 ;
        RECT 97.015 23.055 97.265 23.685 ;
        RECT 96.545 23.515 96.755 24.215 ;
        RECT 96.075 23.135 96.405 23.685 ;
        RECT 94.265 22.765 95.475 23.685 ;
        RECT 94.265 22.225 94.785 23.685 ;
        RECT 94.36 22.225 94.73 24.185 ;
        RECT 88.745 22.745 94.09 23.685 ;
        RECT 92.415 22.745 92.665 24.145 ;
        RECT 91.475 22.745 91.805 24.065 ;
        RECT 88.745 22.225 91.325 23.685 ;
        RECT 88.745 22.225 89.955 24.435 ;
        RECT 88.745 22.225 89.265 24.975 ;
        RECT 88.285 22.79 88.575 24.41 ;
        RECT 84.605 23.515 88.115 24.455 ;
        RECT 87.395 22.905 87.565 24.455 ;
        RECT 86.425 22.985 86.635 24.455 ;
        RECT 84.605 23.515 86.255 24.975 ;
        RECT 84.24 23.015 84.61 23.685 ;
        RECT 83.715 23.515 83.885 24.295 ;
        RECT 82.745 23.515 82.955 24.215 ;
        RECT 82.295 23.055 82.545 23.685 ;
        RECT 81.355 23.135 81.685 23.685 ;
        RECT 80.56 23.515 80.93 24.185 ;
        RECT 79.985 23.135 80.315 23.685 ;
        RECT 74.025 22.745 79.37 23.685 ;
        RECT 78.615 22.745 78.865 24.145 ;
        RECT 77.675 22.745 78.005 24.065 ;
        RECT 75.865 22.745 77.075 24.435 ;
        RECT 74.025 22.225 76.605 23.685 ;
        RECT 75.865 22.225 76.385 24.975 ;
        RECT 74.025 22.225 75.695 24.455 ;
        RECT 74.025 22.225 74.775 24.975 ;
        RECT 73.565 22.79 73.855 24.41 ;
        RECT 72.675 22.905 72.845 23.685 ;
        RECT 71.265 23.515 72.475 24.435 ;
        RECT 71.705 22.985 71.915 24.435 ;
        RECT 71.265 23.515 71.785 24.975 ;
        RECT 70.375 23.515 70.705 24.485 ;
        RECT 69.52 23.015 69.89 23.685 ;
        RECT 69.535 23.015 69.865 24.165 ;
        RECT 68.695 23.515 69.025 24.165 ;
        RECT 67.855 23.515 68.185 24.165 ;
        RECT 67.575 23.055 67.825 23.685 ;
        RECT 67.015 23.515 67.345 24.165 ;
        RECT 66.635 23.135 66.965 23.685 ;
        RECT 66.175 23.515 66.505 24.165 ;
        RECT 64.365 22.745 66.035 23.685 ;
        RECT 62.985 23.515 65.575 24.455 ;
        RECT 64.365 22.225 65.115 24.455 ;
        RECT 62.985 22.745 64.195 24.975 ;
        RECT 61.605 22.745 64.195 23.685 ;
        RECT 59.305 23.515 62.815 24.455 ;
        RECT 61.605 22.225 62.815 24.455 ;
        RECT 60.665 23.135 60.995 24.455 ;
        RECT 59.305 23.515 60.955 24.975 ;
        RECT 58.845 22.79 59.135 24.41 ;
        RECT 57.005 23.515 58.675 24.455 ;
        RECT 57.955 22.905 58.125 24.455 ;
        RECT 57.005 23.515 57.755 24.975 ;
        RECT 56.985 22.985 57.195 23.685 ;
        RECT 56.115 23.515 56.285 24.295 ;
        RECT 55.145 23.515 55.355 24.215 ;
        RECT 54.8 23.015 55.17 23.685 ;
        RECT 52.96 23.515 53.33 24.185 ;
        RECT 52.855 23.055 53.105 23.685 ;
        RECT 51.915 23.135 52.245 23.685 ;
        RECT 49.645 22.745 51.315 23.685 ;
        RECT 51.015 22.745 51.265 24.145 ;
        RECT 50.075 22.745 50.405 24.065 ;
        RECT 49.645 22.225 50.395 23.685 ;
        RECT 48.265 23.515 49.475 24.435 ;
        RECT 48.655 23.035 48.985 24.435 ;
        RECT 48.265 23.515 48.785 24.975 ;
        RECT 44.585 23.515 48.095 24.455 ;
        RECT 46.395 23.035 46.725 24.455 ;
        RECT 44.585 23.515 46.235 24.975 ;
        RECT 44.585 22.765 45.795 24.975 ;
        RECT 44.585 22.225 45.105 24.975 ;
        RECT 44.125 22.79 44.415 24.41 ;
        RECT 42.745 22.765 43.955 24.435 ;
        RECT 42.745 22.225 43.265 24.975 ;
        RECT 40.905 22.745 42.575 24.455 ;
        RECT 40.905 22.225 41.655 24.975 ;
        RECT 35.385 22.745 40.73 24.455 ;
        RECT 35.385 22.225 37.965 24.975 ;
        RECT 29.865 22.745 35.21 24.455 ;
        RECT 29.865 22.225 32.445 24.975 ;
        RECT 29.405 22.79 29.695 24.41 ;
        RECT 26.645 23.515 29.235 24.455 ;
        RECT 28.025 22.765 29.235 24.455 ;
        RECT 28.025 22.225 28.545 24.455 ;
        RECT 26.645 22.745 27.855 24.975 ;
        RECT 26.185 22.225 26.935 23.685 ;
        RECT 25.755 23.515 26.085 24.485 ;
        RECT 20.665 22.745 26.01 23.685 ;
        RECT 24.915 22.745 25.245 24.165 ;
        RECT 24.075 22.745 24.405 24.165 ;
        RECT 23.235 22.745 23.565 24.165 ;
        RECT 20.665 22.225 23.245 23.685 ;
        RECT 22.395 22.225 22.725 24.165 ;
        RECT 21.555 22.225 21.885 24.165 ;
        RECT 19.745 23.515 20.955 24.435 ;
        RECT 15.145 22.745 20.49 23.685 ;
        RECT 19.745 22.745 20.265 24.975 ;
        RECT 17.905 22.745 19.575 24.455 ;
        RECT 17.905 22.745 18.655 24.975 ;
        RECT 15.145 22.745 17.735 24.455 ;
        RECT 15.145 22.225 17.725 24.455 ;
        RECT 15.145 22.225 16.355 24.975 ;
        RECT 14.685 22.79 14.975 24.41 ;
        RECT 13.305 22.765 14.515 24.435 ;
        RECT 13.305 22.225 13.825 24.975 ;
        RECT 10.545 22.745 13.135 24.455 ;
        RECT 10.545 22.225 11.755 24.975 ;
        RECT 10 28.955 189.86 29.125 ;
        RECT 189.025 28.23 189.315 29.85 ;
        RECT 186.265 28.185 188.855 29.895 ;
        RECT 186.265 27.665 187.475 30.415 ;
        RECT 182.585 28.185 186.095 29.895 ;
        RECT 182.585 27.665 184.235 30.415 ;
        RECT 177.065 28.185 182.41 29.895 ;
        RECT 177.065 27.665 179.645 30.415 ;
        RECT 176.605 28.23 176.895 29.85 ;
        RECT 175.225 28.205 176.435 29.875 ;
        RECT 175.225 27.665 175.745 30.415 ;
        RECT 173.385 28.185 175.055 29.895 ;
        RECT 173.385 27.665 174.135 30.415 ;
        RECT 167.865 28.185 173.21 29.895 ;
        RECT 167.865 27.665 170.445 30.415 ;
        RECT 162.345 28.185 167.69 29.895 ;
        RECT 162.345 27.665 164.925 30.415 ;
        RECT 161.885 28.23 162.175 29.85 ;
        RECT 160.505 28.205 161.715 29.875 ;
        RECT 160.505 27.665 161.025 30.415 ;
        RECT 158.665 28.955 160.335 29.895 ;
        RECT 159.515 28.475 159.845 29.895 ;
        RECT 158.665 28.955 159.415 30.415 ;
        RECT 153.145 28.955 158.49 29.895 ;
        RECT 157.255 28.475 157.585 29.895 ;
        RECT 153.145 28.185 156.655 29.895 ;
        RECT 153.145 28.185 155.725 30.415 ;
        RECT 153.145 27.665 154.795 30.415 ;
        RECT 147.625 28.185 152.97 29.895 ;
        RECT 147.625 27.665 150.205 30.415 ;
        RECT 147.165 28.23 147.455 29.85 ;
        RECT 145.325 28.185 146.995 29.125 ;
        RECT 141.645 28.955 146.99 29.895 ;
        RECT 145.325 27.665 146.075 29.895 ;
        RECT 142.565 28.185 145.155 29.895 ;
        RECT 141.645 28.955 144.225 30.415 ;
        RECT 142.565 27.665 143.775 30.415 ;
        RECT 141.675 28.345 141.845 30.415 ;
        RECT 140.715 28.955 141.045 29.605 ;
        RECT 140.705 28.425 140.915 29.125 ;
        RECT 138.52 28.455 138.89 29.125 ;
        RECT 138.455 28.955 138.785 29.605 ;
        RECT 136.585 28.955 137.795 29.875 ;
        RECT 136.585 28.955 137.105 30.415 ;
        RECT 136.575 28.495 136.825 29.125 ;
        RECT 132.905 28.955 136.415 29.895 ;
        RECT 135.635 28.575 135.965 29.895 ;
        RECT 132.905 28.955 134.555 30.415 ;
        RECT 132.905 28.205 134.115 30.415 ;
        RECT 132.905 27.665 133.425 30.415 ;
        RECT 132.445 28.23 132.735 29.85 ;
        RECT 128.765 28.955 132.275 29.895 ;
        RECT 131.095 28.345 131.265 29.895 ;
        RECT 128.765 28.955 130.415 30.415 ;
        RECT 130.125 28.425 130.335 30.415 ;
        RECT 123.245 28.955 128.59 29.895 ;
        RECT 127.94 28.455 128.31 29.895 ;
        RECT 125.995 28.495 126.245 29.895 ;
        RECT 123.245 28.955 125.825 30.415 ;
        RECT 125.055 28.575 125.385 30.415 ;
        RECT 123.245 28.205 124.455 30.415 ;
        RECT 123.245 27.665 123.765 30.415 ;
        RECT 122.255 28.475 122.585 29.605 ;
        RECT 119.995 28.475 120.325 29.605 ;
        RECT 118.185 28.205 119.395 29.875 ;
        RECT 118.185 27.665 118.705 30.415 ;
        RECT 117.725 28.23 118.015 29.85 ;
        RECT 116.345 28.205 117.555 29.875 ;
        RECT 116.345 27.665 116.865 30.415 ;
        RECT 114.505 28.185 116.175 29.895 ;
        RECT 114.505 27.665 115.255 30.415 ;
        RECT 108.985 28.185 114.33 29.895 ;
        RECT 108.985 27.665 111.565 30.415 ;
        RECT 103.465 28.185 108.81 29.895 ;
        RECT 103.465 27.665 106.045 30.415 ;
        RECT 103.005 28.23 103.295 29.85 ;
        RECT 101.625 28.205 102.835 29.125 ;
        RECT 97.485 28.955 102.83 29.895 ;
        RECT 101.625 27.665 102.145 29.895 ;
        RECT 99.785 28.185 101.455 29.895 ;
        RECT 99.785 27.665 100.535 29.895 ;
        RECT 97.485 28.955 100.065 30.415 ;
        RECT 94.265 28.185 99.61 29.125 ;
        RECT 94.265 27.665 96.845 29.125 ;
        RECT 96.495 27.665 96.825 29.605 ;
        RECT 94.235 28.955 94.565 29.605 ;
        RECT 88.745 28.185 94.09 29.125 ;
        RECT 92.425 28.185 93.635 29.875 ;
        RECT 92.425 28.185 92.945 30.415 ;
        RECT 88.745 28.185 92.255 29.895 ;
        RECT 88.745 27.665 91.325 29.895 ;
        RECT 88.745 27.665 90.395 30.415 ;
        RECT 88.285 28.23 88.575 29.85 ;
        RECT 86.905 28.205 88.115 29.875 ;
        RECT 86.905 27.665 87.425 30.415 ;
        RECT 85.065 28.185 86.735 29.895 ;
        RECT 85.065 27.665 85.815 29.895 ;
        RECT 84.145 28.955 85.355 30.415 ;
        RECT 79.545 28.185 84.89 29.125 ;
        RECT 83.155 28.185 83.485 29.605 ;
        RECT 79.545 27.665 82.125 29.125 ;
        RECT 80.895 27.665 81.225 29.605 ;
        RECT 77.705 28.955 80.295 29.895 ;
        RECT 74.025 28.185 79.37 29.125 ;
        RECT 77.705 28.185 78.915 30.415 ;
        RECT 76.715 28.185 77.045 29.605 ;
        RECT 74.025 27.665 76.605 29.125 ;
        RECT 74.455 27.665 74.785 29.605 ;
        RECT 73.565 28.23 73.855 29.85 ;
        RECT 72.185 28.205 73.395 29.875 ;
        RECT 72.185 27.665 72.705 30.415 ;
        RECT 66.665 28.955 72.01 29.895 ;
        RECT 71.255 28.475 71.585 29.895 ;
        RECT 68.995 28.475 69.325 29.895 ;
        RECT 66.665 28.955 69.245 30.415 ;
        RECT 66.665 28.185 68.335 30.415 ;
        RECT 66.665 27.665 67.415 30.415 ;
        RECT 65.775 28.345 65.945 29.735 ;
        RECT 64.805 28.425 65.015 29.655 ;
        RECT 62.62 28.455 62.99 29.625 ;
        RECT 60.675 28.495 60.925 29.585 ;
        RECT 59.735 28.575 60.065 29.505 ;
        RECT 58.845 28.23 59.135 29.85 ;
        RECT 55.165 28.185 58.675 29.895 ;
        RECT 55.165 27.665 56.815 30.415 ;
        RECT 49.645 28.185 54.99 29.895 ;
        RECT 49.645 27.665 52.225 30.415 ;
        RECT 48.655 28.475 48.985 29.605 ;
        RECT 46.395 28.475 46.725 29.605 ;
        RECT 44.585 28.205 45.795 29.875 ;
        RECT 44.585 27.665 45.105 30.415 ;
        RECT 44.125 28.23 44.415 29.85 ;
        RECT 42.745 28.205 43.955 29.875 ;
        RECT 42.745 27.665 43.265 30.415 ;
        RECT 40.905 28.185 42.575 29.895 ;
        RECT 40.905 27.665 41.655 30.415 ;
        RECT 35.385 28.955 40.73 29.895 ;
        RECT 39.975 28.475 40.305 29.895 ;
        RECT 39.135 28.475 39.465 29.895 ;
        RECT 38.295 28.475 38.625 29.895 ;
        RECT 35.385 28.955 37.965 30.415 ;
        RECT 37.455 28.475 37.785 30.415 ;
        RECT 36.615 28.475 36.945 30.415 ;
        RECT 35.775 28.155 36.105 30.415 ;
        RECT 29.865 28.185 35.21 29.895 ;
        RECT 29.865 27.665 32.445 30.415 ;
        RECT 29.405 28.23 29.695 29.85 ;
        RECT 28.025 28.205 29.235 29.875 ;
        RECT 28.025 27.665 28.545 30.415 ;
        RECT 26.185 28.185 27.855 29.895 ;
        RECT 26.185 27.665 26.935 30.415 ;
        RECT 20.665 28.185 26.01 29.895 ;
        RECT 20.665 27.665 23.245 30.415 ;
        RECT 15.145 28.185 20.49 29.895 ;
        RECT 15.145 27.665 17.725 30.415 ;
        RECT 14.685 28.23 14.975 29.85 ;
        RECT 13.305 28.205 14.515 29.875 ;
        RECT 13.305 27.665 13.825 30.415 ;
        RECT 10.545 28.185 13.135 29.895 ;
        RECT 10.545 27.665 11.755 30.415 ;
        RECT 10 34.395 189.86 34.565 ;
        RECT 189.025 33.67 189.315 35.29 ;
        RECT 186.265 33.625 188.855 35.335 ;
        RECT 186.265 33.105 187.475 35.855 ;
        RECT 182.585 33.625 186.095 35.335 ;
        RECT 182.585 33.105 184.235 35.855 ;
        RECT 177.065 33.625 182.41 35.335 ;
        RECT 177.065 33.105 179.645 35.855 ;
        RECT 176.605 33.67 176.895 35.29 ;
        RECT 175.225 33.645 176.435 35.315 ;
        RECT 175.225 33.105 175.745 35.855 ;
        RECT 173.385 33.625 175.055 35.335 ;
        RECT 173.385 33.105 174.135 35.855 ;
        RECT 167.865 33.625 173.21 35.335 ;
        RECT 167.865 33.105 170.445 35.855 ;
        RECT 162.345 33.625 167.69 35.335 ;
        RECT 162.345 33.105 164.925 35.855 ;
        RECT 161.885 33.67 162.175 35.29 ;
        RECT 160.505 33.645 161.715 35.315 ;
        RECT 160.505 33.105 161.025 35.855 ;
        RECT 158.665 33.625 160.335 35.335 ;
        RECT 158.665 33.105 159.415 35.855 ;
        RECT 153.145 33.625 158.49 35.335 ;
        RECT 153.145 33.105 155.725 35.855 ;
        RECT 147.625 33.625 152.97 35.335 ;
        RECT 147.625 33.105 150.205 35.855 ;
        RECT 147.165 33.67 147.455 35.29 ;
        RECT 145.785 33.645 146.995 35.315 ;
        RECT 145.785 33.105 146.305 35.855 ;
        RECT 143.945 33.625 145.615 35.335 ;
        RECT 143.945 33.105 144.695 35.855 ;
        RECT 138.425 33.625 143.77 35.335 ;
        RECT 138.425 33.105 141.005 35.855 ;
        RECT 132.905 33.625 138.25 35.335 ;
        RECT 132.905 33.105 135.485 35.855 ;
        RECT 132.445 33.67 132.735 35.29 ;
        RECT 131.065 33.625 132.275 35.315 ;
        RECT 131.065 33.625 131.585 35.855 ;
        RECT 129.685 33.625 132.275 34.565 ;
        RECT 129.685 33.105 130.895 35.335 ;
        RECT 129.225 34.395 129.975 35.855 ;
        RECT 126.005 33.625 129.515 34.565 ;
        RECT 123.705 34.395 129.05 35.335 ;
        RECT 126.005 33.105 127.655 35.335 ;
        RECT 123.705 34.395 126.285 35.855 ;
        RECT 120.485 33.625 125.83 34.565 ;
        RECT 118.185 34.395 123.53 35.335 ;
        RECT 120.485 33.105 123.065 35.335 ;
        RECT 118.185 34.395 120.765 35.855 ;
        RECT 120.045 33.575 120.275 35.855 ;
        RECT 119.165 33.575 119.375 35.855 ;
        RECT 117.725 33.67 118.015 35.29 ;
        RECT 116.345 33.645 117.555 35.315 ;
        RECT 116.345 33.105 116.865 35.855 ;
        RECT 114.505 33.625 116.175 35.335 ;
        RECT 114.505 33.105 115.255 35.855 ;
        RECT 108.985 33.625 114.33 35.335 ;
        RECT 108.985 33.105 111.565 35.855 ;
        RECT 103.465 33.625 108.81 35.335 ;
        RECT 103.465 33.105 106.045 35.855 ;
        RECT 103.005 33.67 103.295 35.29 ;
        RECT 101.625 33.645 102.835 35.315 ;
        RECT 101.625 33.105 102.145 35.855 ;
        RECT 99.785 33.625 101.455 35.335 ;
        RECT 99.785 33.105 100.535 35.855 ;
        RECT 94.265 33.625 99.61 35.335 ;
        RECT 94.265 33.105 96.845 35.855 ;
        RECT 88.745 33.625 94.09 35.335 ;
        RECT 88.745 33.105 91.325 35.855 ;
        RECT 88.285 33.67 88.575 35.29 ;
        RECT 86.905 33.645 88.115 35.315 ;
        RECT 86.905 33.105 87.425 35.855 ;
        RECT 85.065 33.625 86.735 35.335 ;
        RECT 85.065 33.105 85.815 35.855 ;
      LAYER met1 ;
        RECT 10 12.48 190 12.96 ;
        RECT 10 17.92 190 18.4 ;
        RECT 10 23.36 190 23.84 ;
        RECT 10 28.8 190 29.28 ;
        RECT 10 34.24 190 34.72 ;
        RECT 10 39.68 190 40.16 ;
        RECT 10 45.12 190 45.6 ;
        RECT 10 50.56 190 51.04 ;
        RECT 10 56 190 56.48 ;
      LAYER met4 ;
        RECT 188.23 37.9 189.65 39.9 ;
        RECT 188.23 17.5 189.65 19.5 ;
        RECT 188.47 10 189.41 60 ;
        RECT 182.71 37.9 184.13 39.9 ;
        RECT 182.71 17.5 184.13 19.5 ;
        RECT 182.95 10 183.89 60 ;
        RECT 177.19 37.9 178.61 39.9 ;
        RECT 177.19 17.5 178.61 19.5 ;
        RECT 177.43 10 178.37 60 ;
        RECT 171.67 37.9 173.09 39.9 ;
        RECT 171.67 17.5 173.09 19.5 ;
        RECT 171.91 10 172.85 60 ;
        RECT 166.15 37.9 167.57 39.9 ;
        RECT 166.15 17.5 167.57 19.5 ;
        RECT 166.39 10 167.33 60 ;
        RECT 160.63 37.9 162.05 39.9 ;
        RECT 160.63 17.5 162.05 19.5 ;
        RECT 160.87 10 161.81 60 ;
        RECT 155.11 37.9 156.53 39.9 ;
        RECT 155.11 17.5 156.53 19.5 ;
        RECT 155.35 10 156.29 60 ;
        RECT 149.59 37.9 151.01 39.9 ;
        RECT 149.59 17.5 151.01 19.5 ;
        RECT 149.83 10 150.77 60 ;
        RECT 144.07 37.9 145.49 39.9 ;
        RECT 144.07 17.5 145.49 19.5 ;
        RECT 144.31 10 145.25 60 ;
        RECT 138.55 37.9 139.97 39.9 ;
        RECT 138.55 17.5 139.97 19.5 ;
        RECT 138.79 10 139.73 60 ;
        RECT 133.03 37.9 134.45 39.9 ;
        RECT 133.03 17.5 134.45 19.5 ;
        RECT 133.27 10 134.21 60 ;
        RECT 127.51 37.9 128.93 39.9 ;
        RECT 127.51 17.5 128.93 19.5 ;
        RECT 127.75 10 128.69 60 ;
        RECT 121.99 37.9 123.41 39.9 ;
        RECT 121.99 17.5 123.41 19.5 ;
        RECT 122.23 10 123.17 60 ;
        RECT 116.47 37.9 117.89 39.9 ;
        RECT 116.47 17.5 117.89 19.5 ;
        RECT 116.71 10 117.65 60 ;
        RECT 110.95 37.9 112.37 39.9 ;
        RECT 110.95 17.5 112.37 19.5 ;
        RECT 111.19 10 112.13 60 ;
        RECT 105.43 37.9 106.85 39.9 ;
        RECT 105.43 17.5 106.85 19.5 ;
        RECT 105.67 10 106.61 60 ;
        RECT 99.91 37.9 101.33 39.9 ;
        RECT 99.91 17.5 101.33 19.5 ;
        RECT 100.15 10 101.09 60 ;
        RECT 94.39 37.9 95.81 39.9 ;
        RECT 94.39 17.5 95.81 19.5 ;
        RECT 94.63 10 95.57 60 ;
        RECT 88.87 37.9 90.29 39.9 ;
        RECT 88.87 17.5 90.29 19.5 ;
        RECT 89.11 10 90.05 60 ;
        RECT 83.35 37.9 84.77 39.9 ;
        RECT 83.35 17.5 84.77 19.5 ;
        RECT 83.59 10 84.53 60 ;
        RECT 77.83 37.9 79.25 39.9 ;
        RECT 77.83 17.5 79.25 19.5 ;
        RECT 78.07 10 79.01 60 ;
        RECT 72.31 37.9 73.73 39.9 ;
        RECT 72.31 17.5 73.73 19.5 ;
        RECT 72.55 10 73.49 60 ;
        RECT 66.79 37.9 68.21 39.9 ;
        RECT 66.79 17.5 68.21 19.5 ;
        RECT 67.03 10 67.97 60 ;
        RECT 61.27 37.9 62.69 39.9 ;
        RECT 61.27 17.5 62.69 19.5 ;
        RECT 61.51 10 62.45 60 ;
        RECT 55.75 37.9 57.17 39.9 ;
        RECT 55.75 17.5 57.17 19.5 ;
        RECT 55.99 10 56.93 60 ;
        RECT 50.23 37.9 51.65 39.9 ;
        RECT 50.23 17.5 51.65 19.5 ;
        RECT 50.47 10 51.41 60 ;
        RECT 44.71 37.9 46.13 39.9 ;
        RECT 44.71 17.5 46.13 19.5 ;
        RECT 44.95 10 45.89 60 ;
        RECT 39.19 37.9 40.61 39.9 ;
        RECT 39.19 17.5 40.61 19.5 ;
        RECT 39.43 10 40.37 60 ;
        RECT 33.67 37.9 35.09 39.9 ;
        RECT 33.67 17.5 35.09 19.5 ;
        RECT 33.91 10 34.85 60 ;
        RECT 28.15 37.9 29.57 39.9 ;
        RECT 28.15 17.5 29.57 19.5 ;
        RECT 28.39 10 29.33 60 ;
        RECT 22.63 37.9 24.05 39.9 ;
        RECT 22.63 17.5 24.05 19.5 ;
        RECT 22.87 10 23.81 60 ;
        RECT 17.11 37.9 18.53 39.9 ;
        RECT 17.11 17.5 18.53 19.5 ;
        RECT 17.35 10 18.29 60 ;
        RECT 11.59 37.9 13.01 39.9 ;
        RECT 11.59 17.5 13.01 19.5 ;
        RECT 11.83 10 12.77 60 ;
      LAYER met3 ;
        RECT 10 11.47 190 11.93 ;
        RECT 10 15.55 190 16.01 ;
        RECT 10 19.63 190 20.09 ;
        RECT 10 23.71 190 24.17 ;
        RECT 10 27.79 190 28.25 ;
        RECT 10 31.87 190 32.33 ;
        RECT 10 35.95 190 36.41 ;
        RECT 10 40.03 190 40.49 ;
        RECT 10 44.11 190 44.57 ;
        RECT 10 48.19 190 48.65 ;
        RECT 10 52.27 190 52.73 ;
        RECT 10 56.35 190 56.81 ;
      LAYER met2 ;
        RECT 187.54 10 188.04 60 ;
        RECT 184.78 10 185.28 60 ;
        RECT 182.02 10 182.52 60 ;
        RECT 179.26 10 179.76 60 ;
        RECT 176.5 10 177 60 ;
        RECT 173.74 10 174.24 60 ;
        RECT 170.98 10 171.48 60 ;
        RECT 168.22 10 168.72 60 ;
        RECT 165.46 10 165.96 60 ;
        RECT 162.7 10 163.2 60 ;
        RECT 159.94 10 160.44 60 ;
        RECT 157.18 10 157.68 60 ;
        RECT 154.42 10 154.92 60 ;
        RECT 151.66 10 152.16 60 ;
        RECT 148.9 10 149.4 60 ;
        RECT 146.14 10 146.64 60 ;
        RECT 143.38 10 143.88 60 ;
        RECT 140.62 10 141.12 60 ;
        RECT 137.86 10 138.36 60 ;
        RECT 135.1 10 135.6 60 ;
        RECT 132.34 10 132.84 60 ;
        RECT 129.58 10 130.08 60 ;
        RECT 126.82 10 127.32 60 ;
        RECT 124.06 10 124.56 60 ;
        RECT 121.3 10 121.8 60 ;
        RECT 118.54 10 119.04 60 ;
        RECT 115.78 10 116.28 60 ;
        RECT 113.02 10 113.52 60 ;
        RECT 110.26 10 110.76 60 ;
        RECT 107.5 10 108 60 ;
        RECT 104.74 10 105.24 60 ;
        RECT 101.98 10 102.48 60 ;
        RECT 99.22 10 99.72 60 ;
        RECT 96.46 10 96.96 60 ;
        RECT 93.7 10 94.2 60 ;
        RECT 90.94 10 91.44 60 ;
        RECT 88.18 10 88.68 60 ;
        RECT 85.42 10 85.92 60 ;
        RECT 82.66 10 83.16 60 ;
        RECT 79.9 10 80.4 60 ;
        RECT 77.14 10 77.64 60 ;
        RECT 74.38 10 74.88 60 ;
        RECT 71.62 10 72.12 60 ;
        RECT 68.86 10 69.36 60 ;
        RECT 66.1 10 66.6 60 ;
        RECT 63.34 10 63.84 60 ;
        RECT 60.58 10 61.08 60 ;
        RECT 57.82 10 58.32 60 ;
        RECT 55.06 10 55.56 60 ;
        RECT 52.3 10 52.8 60 ;
        RECT 49.54 10 50.04 60 ;
        RECT 46.78 10 47.28 60 ;
        RECT 44.02 10 44.52 60 ;
        RECT 41.26 10 41.76 60 ;
        RECT 38.5 10 39 60 ;
        RECT 35.74 10 36.24 60 ;
        RECT 32.98 10 33.48 60 ;
        RECT 30.22 10 30.72 60 ;
        RECT 27.46 10 27.96 60 ;
        RECT 24.7 10 25.2 60 ;
        RECT 21.94 10 22.44 60 ;
        RECT 19.18 10 19.68 60 ;
        RECT 16.42 10 16.92 60 ;
        RECT 13.66 10 14.16 60 ;
        RECT 10.9 10 11.4 60 ;
      LAYER via3 ;
        RECT 12 56.48 12.2 56.68 ;
        RECT 12 52.4 12.2 52.6 ;
        RECT 12 48.32 12.2 48.52 ;
        RECT 12 44.24 12.2 44.44 ;
        RECT 12 40.16 12.2 40.36 ;
        RECT 12 36.08 12.2 36.28 ;
        RECT 12 32 12.2 32.2 ;
        RECT 12 27.92 12.2 28.12 ;
        RECT 12 23.84 12.2 24.04 ;
        RECT 12 19.76 12.2 19.96 ;
        RECT 12 15.68 12.2 15.88 ;
        RECT 12 11.6 12.2 11.8 ;
        RECT 12.4 56.48 12.6 56.68 ;
        RECT 12.4 52.4 12.6 52.6 ;
        RECT 12.4 48.32 12.6 48.52 ;
        RECT 12.4 44.24 12.6 44.44 ;
        RECT 12.4 40.16 12.6 40.36 ;
        RECT 12.4 36.08 12.6 36.28 ;
        RECT 12.4 32 12.6 32.2 ;
        RECT 12.4 27.92 12.6 28.12 ;
        RECT 12.4 23.84 12.6 24.04 ;
        RECT 12.4 19.76 12.6 19.96 ;
        RECT 12.4 15.68 12.6 15.88 ;
        RECT 12.4 11.6 12.6 11.8 ;
        RECT 17.52 56.48 17.72 56.68 ;
        RECT 17.52 52.4 17.72 52.6 ;
        RECT 17.52 48.32 17.72 48.52 ;
        RECT 17.52 44.24 17.72 44.44 ;
        RECT 17.52 40.16 17.72 40.36 ;
        RECT 17.52 36.08 17.72 36.28 ;
        RECT 17.52 32 17.72 32.2 ;
        RECT 17.52 27.92 17.72 28.12 ;
        RECT 17.52 23.84 17.72 24.04 ;
        RECT 17.52 19.76 17.72 19.96 ;
        RECT 17.52 15.68 17.72 15.88 ;
        RECT 17.52 11.6 17.72 11.8 ;
        RECT 17.92 56.48 18.12 56.68 ;
        RECT 17.92 52.4 18.12 52.6 ;
        RECT 17.92 48.32 18.12 48.52 ;
        RECT 17.92 44.24 18.12 44.44 ;
        RECT 17.92 40.16 18.12 40.36 ;
        RECT 17.92 36.08 18.12 36.28 ;
        RECT 17.92 32 18.12 32.2 ;
        RECT 17.92 27.92 18.12 28.12 ;
        RECT 17.92 23.84 18.12 24.04 ;
        RECT 17.92 19.76 18.12 19.96 ;
        RECT 17.92 15.68 18.12 15.88 ;
        RECT 17.92 11.6 18.12 11.8 ;
        RECT 23.04 56.48 23.24 56.68 ;
        RECT 23.04 52.4 23.24 52.6 ;
        RECT 23.04 48.32 23.24 48.52 ;
        RECT 23.04 44.24 23.24 44.44 ;
        RECT 23.04 40.16 23.24 40.36 ;
        RECT 23.04 36.08 23.24 36.28 ;
        RECT 23.04 32 23.24 32.2 ;
        RECT 23.04 27.92 23.24 28.12 ;
        RECT 23.04 23.84 23.24 24.04 ;
        RECT 23.04 19.76 23.24 19.96 ;
        RECT 23.04 15.68 23.24 15.88 ;
        RECT 23.04 11.6 23.24 11.8 ;
        RECT 23.44 56.48 23.64 56.68 ;
        RECT 23.44 52.4 23.64 52.6 ;
        RECT 23.44 48.32 23.64 48.52 ;
        RECT 23.44 44.24 23.64 44.44 ;
        RECT 23.44 40.16 23.64 40.36 ;
        RECT 23.44 36.08 23.64 36.28 ;
        RECT 23.44 32 23.64 32.2 ;
        RECT 23.44 27.92 23.64 28.12 ;
        RECT 23.44 23.84 23.64 24.04 ;
        RECT 23.44 19.76 23.64 19.96 ;
        RECT 23.44 15.68 23.64 15.88 ;
        RECT 23.44 11.6 23.64 11.8 ;
        RECT 28.56 56.48 28.76 56.68 ;
        RECT 28.56 52.4 28.76 52.6 ;
        RECT 28.56 48.32 28.76 48.52 ;
        RECT 28.56 44.24 28.76 44.44 ;
        RECT 28.56 40.16 28.76 40.36 ;
        RECT 28.56 36.08 28.76 36.28 ;
        RECT 28.56 32 28.76 32.2 ;
        RECT 28.56 27.92 28.76 28.12 ;
        RECT 28.56 23.84 28.76 24.04 ;
        RECT 28.56 19.76 28.76 19.96 ;
        RECT 28.56 15.68 28.76 15.88 ;
        RECT 28.56 11.6 28.76 11.8 ;
        RECT 28.96 56.48 29.16 56.68 ;
        RECT 28.96 52.4 29.16 52.6 ;
        RECT 28.96 48.32 29.16 48.52 ;
        RECT 28.96 44.24 29.16 44.44 ;
        RECT 28.96 40.16 29.16 40.36 ;
        RECT 28.96 36.08 29.16 36.28 ;
        RECT 28.96 32 29.16 32.2 ;
        RECT 28.96 27.92 29.16 28.12 ;
        RECT 28.96 23.84 29.16 24.04 ;
        RECT 28.96 19.76 29.16 19.96 ;
        RECT 28.96 15.68 29.16 15.88 ;
        RECT 28.96 11.6 29.16 11.8 ;
        RECT 34.08 56.48 34.28 56.68 ;
        RECT 34.08 52.4 34.28 52.6 ;
        RECT 34.08 48.32 34.28 48.52 ;
        RECT 34.08 44.24 34.28 44.44 ;
        RECT 34.08 40.16 34.28 40.36 ;
        RECT 34.08 36.08 34.28 36.28 ;
        RECT 34.08 32 34.28 32.2 ;
        RECT 34.08 27.92 34.28 28.12 ;
        RECT 34.08 23.84 34.28 24.04 ;
        RECT 34.08 19.76 34.28 19.96 ;
        RECT 34.08 15.68 34.28 15.88 ;
        RECT 34.08 11.6 34.28 11.8 ;
        RECT 34.48 56.48 34.68 56.68 ;
        RECT 34.48 52.4 34.68 52.6 ;
        RECT 34.48 48.32 34.68 48.52 ;
        RECT 34.48 44.24 34.68 44.44 ;
        RECT 34.48 40.16 34.68 40.36 ;
        RECT 34.48 36.08 34.68 36.28 ;
        RECT 34.48 32 34.68 32.2 ;
        RECT 34.48 27.92 34.68 28.12 ;
        RECT 34.48 23.84 34.68 24.04 ;
        RECT 34.48 19.76 34.68 19.96 ;
        RECT 34.48 15.68 34.68 15.88 ;
        RECT 34.48 11.6 34.68 11.8 ;
        RECT 39.6 56.48 39.8 56.68 ;
        RECT 39.6 52.4 39.8 52.6 ;
        RECT 39.6 48.32 39.8 48.52 ;
        RECT 39.6 44.24 39.8 44.44 ;
        RECT 39.6 40.16 39.8 40.36 ;
        RECT 39.6 36.08 39.8 36.28 ;
        RECT 39.6 32 39.8 32.2 ;
        RECT 39.6 27.92 39.8 28.12 ;
        RECT 39.6 23.84 39.8 24.04 ;
        RECT 39.6 19.76 39.8 19.96 ;
        RECT 39.6 15.68 39.8 15.88 ;
        RECT 39.6 11.6 39.8 11.8 ;
        RECT 40 56.48 40.2 56.68 ;
        RECT 40 52.4 40.2 52.6 ;
        RECT 40 48.32 40.2 48.52 ;
        RECT 40 44.24 40.2 44.44 ;
        RECT 40 40.16 40.2 40.36 ;
        RECT 40 36.08 40.2 36.28 ;
        RECT 40 32 40.2 32.2 ;
        RECT 40 27.92 40.2 28.12 ;
        RECT 40 23.84 40.2 24.04 ;
        RECT 40 19.76 40.2 19.96 ;
        RECT 40 15.68 40.2 15.88 ;
        RECT 40 11.6 40.2 11.8 ;
        RECT 45.12 56.48 45.32 56.68 ;
        RECT 45.12 52.4 45.32 52.6 ;
        RECT 45.12 48.32 45.32 48.52 ;
        RECT 45.12 44.24 45.32 44.44 ;
        RECT 45.12 40.16 45.32 40.36 ;
        RECT 45.12 36.08 45.32 36.28 ;
        RECT 45.12 32 45.32 32.2 ;
        RECT 45.12 27.92 45.32 28.12 ;
        RECT 45.12 23.84 45.32 24.04 ;
        RECT 45.12 19.76 45.32 19.96 ;
        RECT 45.12 15.68 45.32 15.88 ;
        RECT 45.12 11.6 45.32 11.8 ;
        RECT 45.52 56.48 45.72 56.68 ;
        RECT 45.52 52.4 45.72 52.6 ;
        RECT 45.52 48.32 45.72 48.52 ;
        RECT 45.52 44.24 45.72 44.44 ;
        RECT 45.52 40.16 45.72 40.36 ;
        RECT 45.52 36.08 45.72 36.28 ;
        RECT 45.52 32 45.72 32.2 ;
        RECT 45.52 27.92 45.72 28.12 ;
        RECT 45.52 23.84 45.72 24.04 ;
        RECT 45.52 19.76 45.72 19.96 ;
        RECT 45.52 15.68 45.72 15.88 ;
        RECT 45.52 11.6 45.72 11.8 ;
        RECT 50.64 56.48 50.84 56.68 ;
        RECT 50.64 52.4 50.84 52.6 ;
        RECT 50.64 48.32 50.84 48.52 ;
        RECT 50.64 44.24 50.84 44.44 ;
        RECT 50.64 40.16 50.84 40.36 ;
        RECT 50.64 36.08 50.84 36.28 ;
        RECT 50.64 32 50.84 32.2 ;
        RECT 50.64 27.92 50.84 28.12 ;
        RECT 50.64 23.84 50.84 24.04 ;
        RECT 50.64 19.76 50.84 19.96 ;
        RECT 50.64 15.68 50.84 15.88 ;
        RECT 50.64 11.6 50.84 11.8 ;
        RECT 51.04 56.48 51.24 56.68 ;
        RECT 51.04 52.4 51.24 52.6 ;
        RECT 51.04 48.32 51.24 48.52 ;
        RECT 51.04 44.24 51.24 44.44 ;
        RECT 51.04 40.16 51.24 40.36 ;
        RECT 51.04 36.08 51.24 36.28 ;
        RECT 51.04 32 51.24 32.2 ;
        RECT 51.04 27.92 51.24 28.12 ;
        RECT 51.04 23.84 51.24 24.04 ;
        RECT 51.04 19.76 51.24 19.96 ;
        RECT 51.04 15.68 51.24 15.88 ;
        RECT 51.04 11.6 51.24 11.8 ;
        RECT 56.16 56.48 56.36 56.68 ;
        RECT 56.16 52.4 56.36 52.6 ;
        RECT 56.16 48.32 56.36 48.52 ;
        RECT 56.16 44.24 56.36 44.44 ;
        RECT 56.16 40.16 56.36 40.36 ;
        RECT 56.16 36.08 56.36 36.28 ;
        RECT 56.16 32 56.36 32.2 ;
        RECT 56.16 27.92 56.36 28.12 ;
        RECT 56.16 23.84 56.36 24.04 ;
        RECT 56.16 19.76 56.36 19.96 ;
        RECT 56.16 15.68 56.36 15.88 ;
        RECT 56.16 11.6 56.36 11.8 ;
        RECT 56.56 56.48 56.76 56.68 ;
        RECT 56.56 52.4 56.76 52.6 ;
        RECT 56.56 48.32 56.76 48.52 ;
        RECT 56.56 44.24 56.76 44.44 ;
        RECT 56.56 40.16 56.76 40.36 ;
        RECT 56.56 36.08 56.76 36.28 ;
        RECT 56.56 32 56.76 32.2 ;
        RECT 56.56 27.92 56.76 28.12 ;
        RECT 56.56 23.84 56.76 24.04 ;
        RECT 56.56 19.76 56.76 19.96 ;
        RECT 56.56 15.68 56.76 15.88 ;
        RECT 56.56 11.6 56.76 11.8 ;
        RECT 61.68 56.48 61.88 56.68 ;
        RECT 61.68 52.4 61.88 52.6 ;
        RECT 61.68 48.32 61.88 48.52 ;
        RECT 61.68 44.24 61.88 44.44 ;
        RECT 61.68 40.16 61.88 40.36 ;
        RECT 61.68 36.08 61.88 36.28 ;
        RECT 61.68 32 61.88 32.2 ;
        RECT 61.68 27.92 61.88 28.12 ;
        RECT 61.68 23.84 61.88 24.04 ;
        RECT 61.68 19.76 61.88 19.96 ;
        RECT 61.68 15.68 61.88 15.88 ;
        RECT 61.68 11.6 61.88 11.8 ;
        RECT 62.08 56.48 62.28 56.68 ;
        RECT 62.08 52.4 62.28 52.6 ;
        RECT 62.08 48.32 62.28 48.52 ;
        RECT 62.08 44.24 62.28 44.44 ;
        RECT 62.08 40.16 62.28 40.36 ;
        RECT 62.08 36.08 62.28 36.28 ;
        RECT 62.08 32 62.28 32.2 ;
        RECT 62.08 27.92 62.28 28.12 ;
        RECT 62.08 23.84 62.28 24.04 ;
        RECT 62.08 19.76 62.28 19.96 ;
        RECT 62.08 15.68 62.28 15.88 ;
        RECT 62.08 11.6 62.28 11.8 ;
        RECT 67.2 56.48 67.4 56.68 ;
        RECT 67.2 52.4 67.4 52.6 ;
        RECT 67.2 48.32 67.4 48.52 ;
        RECT 67.2 44.24 67.4 44.44 ;
        RECT 67.2 40.16 67.4 40.36 ;
        RECT 67.2 36.08 67.4 36.28 ;
        RECT 67.2 32 67.4 32.2 ;
        RECT 67.2 27.92 67.4 28.12 ;
        RECT 67.2 23.84 67.4 24.04 ;
        RECT 67.2 19.76 67.4 19.96 ;
        RECT 67.2 15.68 67.4 15.88 ;
        RECT 67.2 11.6 67.4 11.8 ;
        RECT 67.6 56.48 67.8 56.68 ;
        RECT 67.6 52.4 67.8 52.6 ;
        RECT 67.6 48.32 67.8 48.52 ;
        RECT 67.6 44.24 67.8 44.44 ;
        RECT 67.6 40.16 67.8 40.36 ;
        RECT 67.6 36.08 67.8 36.28 ;
        RECT 67.6 32 67.8 32.2 ;
        RECT 67.6 27.92 67.8 28.12 ;
        RECT 67.6 23.84 67.8 24.04 ;
        RECT 67.6 19.76 67.8 19.96 ;
        RECT 67.6 15.68 67.8 15.88 ;
        RECT 67.6 11.6 67.8 11.8 ;
        RECT 72.72 56.48 72.92 56.68 ;
        RECT 72.72 52.4 72.92 52.6 ;
        RECT 72.72 48.32 72.92 48.52 ;
        RECT 72.72 44.24 72.92 44.44 ;
        RECT 72.72 40.16 72.92 40.36 ;
        RECT 72.72 36.08 72.92 36.28 ;
        RECT 72.72 32 72.92 32.2 ;
        RECT 72.72 27.92 72.92 28.12 ;
        RECT 72.72 23.84 72.92 24.04 ;
        RECT 72.72 19.76 72.92 19.96 ;
        RECT 72.72 15.68 72.92 15.88 ;
        RECT 72.72 11.6 72.92 11.8 ;
        RECT 73.12 56.48 73.32 56.68 ;
        RECT 73.12 52.4 73.32 52.6 ;
        RECT 73.12 48.32 73.32 48.52 ;
        RECT 73.12 44.24 73.32 44.44 ;
        RECT 73.12 40.16 73.32 40.36 ;
        RECT 73.12 36.08 73.32 36.28 ;
        RECT 73.12 32 73.32 32.2 ;
        RECT 73.12 27.92 73.32 28.12 ;
        RECT 73.12 23.84 73.32 24.04 ;
        RECT 73.12 19.76 73.32 19.96 ;
        RECT 73.12 15.68 73.32 15.88 ;
        RECT 73.12 11.6 73.32 11.8 ;
        RECT 78.24 56.48 78.44 56.68 ;
        RECT 78.24 52.4 78.44 52.6 ;
        RECT 78.24 48.32 78.44 48.52 ;
        RECT 78.24 44.24 78.44 44.44 ;
        RECT 78.24 40.16 78.44 40.36 ;
        RECT 78.24 36.08 78.44 36.28 ;
        RECT 78.24 32 78.44 32.2 ;
        RECT 78.24 27.92 78.44 28.12 ;
        RECT 78.24 23.84 78.44 24.04 ;
        RECT 78.24 19.76 78.44 19.96 ;
        RECT 78.24 15.68 78.44 15.88 ;
        RECT 78.24 11.6 78.44 11.8 ;
        RECT 78.64 56.48 78.84 56.68 ;
        RECT 78.64 52.4 78.84 52.6 ;
        RECT 78.64 48.32 78.84 48.52 ;
        RECT 78.64 44.24 78.84 44.44 ;
        RECT 78.64 40.16 78.84 40.36 ;
        RECT 78.64 36.08 78.84 36.28 ;
        RECT 78.64 32 78.84 32.2 ;
        RECT 78.64 27.92 78.84 28.12 ;
        RECT 78.64 23.84 78.84 24.04 ;
        RECT 78.64 19.76 78.84 19.96 ;
        RECT 78.64 15.68 78.84 15.88 ;
        RECT 78.64 11.6 78.84 11.8 ;
        RECT 83.76 56.48 83.96 56.68 ;
        RECT 83.76 52.4 83.96 52.6 ;
        RECT 83.76 48.32 83.96 48.52 ;
        RECT 83.76 44.24 83.96 44.44 ;
        RECT 83.76 40.16 83.96 40.36 ;
        RECT 83.76 36.08 83.96 36.28 ;
        RECT 83.76 32 83.96 32.2 ;
        RECT 83.76 27.92 83.96 28.12 ;
        RECT 83.76 23.84 83.96 24.04 ;
        RECT 83.76 19.76 83.96 19.96 ;
        RECT 83.76 15.68 83.96 15.88 ;
        RECT 83.76 11.6 83.96 11.8 ;
        RECT 84.16 56.48 84.36 56.68 ;
        RECT 84.16 52.4 84.36 52.6 ;
        RECT 84.16 48.32 84.36 48.52 ;
        RECT 84.16 44.24 84.36 44.44 ;
        RECT 84.16 40.16 84.36 40.36 ;
        RECT 84.16 36.08 84.36 36.28 ;
        RECT 84.16 32 84.36 32.2 ;
        RECT 84.16 27.92 84.36 28.12 ;
        RECT 84.16 23.84 84.36 24.04 ;
        RECT 84.16 19.76 84.36 19.96 ;
        RECT 84.16 15.68 84.36 15.88 ;
        RECT 84.16 11.6 84.36 11.8 ;
        RECT 89.28 56.48 89.48 56.68 ;
        RECT 89.28 52.4 89.48 52.6 ;
        RECT 89.28 48.32 89.48 48.52 ;
        RECT 89.28 44.24 89.48 44.44 ;
        RECT 89.28 40.16 89.48 40.36 ;
        RECT 89.28 36.08 89.48 36.28 ;
        RECT 89.28 32 89.48 32.2 ;
        RECT 89.28 27.92 89.48 28.12 ;
        RECT 89.28 23.84 89.48 24.04 ;
        RECT 89.28 19.76 89.48 19.96 ;
        RECT 89.28 15.68 89.48 15.88 ;
        RECT 89.28 11.6 89.48 11.8 ;
        RECT 89.68 56.48 89.88 56.68 ;
        RECT 89.68 52.4 89.88 52.6 ;
        RECT 89.68 48.32 89.88 48.52 ;
        RECT 89.68 44.24 89.88 44.44 ;
        RECT 89.68 40.16 89.88 40.36 ;
        RECT 89.68 36.08 89.88 36.28 ;
        RECT 89.68 32 89.88 32.2 ;
        RECT 89.68 27.92 89.88 28.12 ;
        RECT 89.68 23.84 89.88 24.04 ;
        RECT 89.68 19.76 89.88 19.96 ;
        RECT 89.68 15.68 89.88 15.88 ;
        RECT 89.68 11.6 89.88 11.8 ;
        RECT 94.8 56.48 95 56.68 ;
        RECT 94.8 52.4 95 52.6 ;
        RECT 94.8 48.32 95 48.52 ;
        RECT 94.8 44.24 95 44.44 ;
        RECT 94.8 40.16 95 40.36 ;
        RECT 94.8 36.08 95 36.28 ;
        RECT 94.8 32 95 32.2 ;
        RECT 94.8 27.92 95 28.12 ;
        RECT 94.8 23.84 95 24.04 ;
        RECT 94.8 19.76 95 19.96 ;
        RECT 94.8 15.68 95 15.88 ;
        RECT 94.8 11.6 95 11.8 ;
        RECT 95.2 56.48 95.4 56.68 ;
        RECT 95.2 52.4 95.4 52.6 ;
        RECT 95.2 48.32 95.4 48.52 ;
        RECT 95.2 44.24 95.4 44.44 ;
        RECT 95.2 40.16 95.4 40.36 ;
        RECT 95.2 36.08 95.4 36.28 ;
        RECT 95.2 32 95.4 32.2 ;
        RECT 95.2 27.92 95.4 28.12 ;
        RECT 95.2 23.84 95.4 24.04 ;
        RECT 95.2 19.76 95.4 19.96 ;
        RECT 95.2 15.68 95.4 15.88 ;
        RECT 95.2 11.6 95.4 11.8 ;
        RECT 100.32 56.48 100.52 56.68 ;
        RECT 100.32 52.4 100.52 52.6 ;
        RECT 100.32 48.32 100.52 48.52 ;
        RECT 100.32 44.24 100.52 44.44 ;
        RECT 100.32 40.16 100.52 40.36 ;
        RECT 100.32 36.08 100.52 36.28 ;
        RECT 100.32 32 100.52 32.2 ;
        RECT 100.32 27.92 100.52 28.12 ;
        RECT 100.32 23.84 100.52 24.04 ;
        RECT 100.32 19.76 100.52 19.96 ;
        RECT 100.32 15.68 100.52 15.88 ;
        RECT 100.32 11.6 100.52 11.8 ;
        RECT 100.72 56.48 100.92 56.68 ;
        RECT 100.72 52.4 100.92 52.6 ;
        RECT 100.72 48.32 100.92 48.52 ;
        RECT 100.72 44.24 100.92 44.44 ;
        RECT 100.72 40.16 100.92 40.36 ;
        RECT 100.72 36.08 100.92 36.28 ;
        RECT 100.72 32 100.92 32.2 ;
        RECT 100.72 27.92 100.92 28.12 ;
        RECT 100.72 23.84 100.92 24.04 ;
        RECT 100.72 19.76 100.92 19.96 ;
        RECT 100.72 15.68 100.92 15.88 ;
        RECT 100.72 11.6 100.92 11.8 ;
        RECT 105.84 56.48 106.04 56.68 ;
        RECT 105.84 52.4 106.04 52.6 ;
        RECT 105.84 48.32 106.04 48.52 ;
        RECT 105.84 44.24 106.04 44.44 ;
        RECT 105.84 40.16 106.04 40.36 ;
        RECT 105.84 36.08 106.04 36.28 ;
        RECT 105.84 32 106.04 32.2 ;
        RECT 105.84 27.92 106.04 28.12 ;
        RECT 105.84 23.84 106.04 24.04 ;
        RECT 105.84 19.76 106.04 19.96 ;
        RECT 105.84 15.68 106.04 15.88 ;
        RECT 105.84 11.6 106.04 11.8 ;
        RECT 106.24 56.48 106.44 56.68 ;
        RECT 106.24 52.4 106.44 52.6 ;
        RECT 106.24 48.32 106.44 48.52 ;
        RECT 106.24 44.24 106.44 44.44 ;
        RECT 106.24 40.16 106.44 40.36 ;
        RECT 106.24 36.08 106.44 36.28 ;
        RECT 106.24 32 106.44 32.2 ;
        RECT 106.24 27.92 106.44 28.12 ;
        RECT 106.24 23.84 106.44 24.04 ;
        RECT 106.24 19.76 106.44 19.96 ;
        RECT 106.24 15.68 106.44 15.88 ;
        RECT 106.24 11.6 106.44 11.8 ;
        RECT 111.36 56.48 111.56 56.68 ;
        RECT 111.36 52.4 111.56 52.6 ;
        RECT 111.36 48.32 111.56 48.52 ;
        RECT 111.36 44.24 111.56 44.44 ;
        RECT 111.36 40.16 111.56 40.36 ;
        RECT 111.36 36.08 111.56 36.28 ;
        RECT 111.36 32 111.56 32.2 ;
        RECT 111.36 27.92 111.56 28.12 ;
        RECT 111.36 23.84 111.56 24.04 ;
        RECT 111.36 19.76 111.56 19.96 ;
        RECT 111.36 15.68 111.56 15.88 ;
        RECT 111.36 11.6 111.56 11.8 ;
        RECT 111.76 56.48 111.96 56.68 ;
        RECT 111.76 52.4 111.96 52.6 ;
        RECT 111.76 48.32 111.96 48.52 ;
        RECT 111.76 44.24 111.96 44.44 ;
        RECT 111.76 40.16 111.96 40.36 ;
        RECT 111.76 36.08 111.96 36.28 ;
        RECT 111.76 32 111.96 32.2 ;
        RECT 111.76 27.92 111.96 28.12 ;
        RECT 111.76 23.84 111.96 24.04 ;
        RECT 111.76 19.76 111.96 19.96 ;
        RECT 111.76 15.68 111.96 15.88 ;
        RECT 111.76 11.6 111.96 11.8 ;
        RECT 116.88 56.48 117.08 56.68 ;
        RECT 116.88 52.4 117.08 52.6 ;
        RECT 116.88 48.32 117.08 48.52 ;
        RECT 116.88 44.24 117.08 44.44 ;
        RECT 116.88 40.16 117.08 40.36 ;
        RECT 116.88 36.08 117.08 36.28 ;
        RECT 116.88 32 117.08 32.2 ;
        RECT 116.88 27.92 117.08 28.12 ;
        RECT 116.88 23.84 117.08 24.04 ;
        RECT 116.88 19.76 117.08 19.96 ;
        RECT 116.88 15.68 117.08 15.88 ;
        RECT 116.88 11.6 117.08 11.8 ;
        RECT 117.28 56.48 117.48 56.68 ;
        RECT 117.28 52.4 117.48 52.6 ;
        RECT 117.28 48.32 117.48 48.52 ;
        RECT 117.28 44.24 117.48 44.44 ;
        RECT 117.28 40.16 117.48 40.36 ;
        RECT 117.28 36.08 117.48 36.28 ;
        RECT 117.28 32 117.48 32.2 ;
        RECT 117.28 27.92 117.48 28.12 ;
        RECT 117.28 23.84 117.48 24.04 ;
        RECT 117.28 19.76 117.48 19.96 ;
        RECT 117.28 15.68 117.48 15.88 ;
        RECT 117.28 11.6 117.48 11.8 ;
        RECT 122.4 56.48 122.6 56.68 ;
        RECT 122.4 52.4 122.6 52.6 ;
        RECT 122.4 48.32 122.6 48.52 ;
        RECT 122.4 44.24 122.6 44.44 ;
        RECT 122.4 40.16 122.6 40.36 ;
        RECT 122.4 36.08 122.6 36.28 ;
        RECT 122.4 32 122.6 32.2 ;
        RECT 122.4 27.92 122.6 28.12 ;
        RECT 122.4 23.84 122.6 24.04 ;
        RECT 122.4 19.76 122.6 19.96 ;
        RECT 122.4 15.68 122.6 15.88 ;
        RECT 122.4 11.6 122.6 11.8 ;
        RECT 122.8 56.48 123 56.68 ;
        RECT 122.8 52.4 123 52.6 ;
        RECT 122.8 48.32 123 48.52 ;
        RECT 122.8 44.24 123 44.44 ;
        RECT 122.8 40.16 123 40.36 ;
        RECT 122.8 36.08 123 36.28 ;
        RECT 122.8 32 123 32.2 ;
        RECT 122.8 27.92 123 28.12 ;
        RECT 122.8 23.84 123 24.04 ;
        RECT 122.8 19.76 123 19.96 ;
        RECT 122.8 15.68 123 15.88 ;
        RECT 122.8 11.6 123 11.8 ;
        RECT 127.92 56.48 128.12 56.68 ;
        RECT 127.92 52.4 128.12 52.6 ;
        RECT 127.92 48.32 128.12 48.52 ;
        RECT 127.92 44.24 128.12 44.44 ;
        RECT 127.92 40.16 128.12 40.36 ;
        RECT 127.92 36.08 128.12 36.28 ;
        RECT 127.92 32 128.12 32.2 ;
        RECT 127.92 27.92 128.12 28.12 ;
        RECT 127.92 23.84 128.12 24.04 ;
        RECT 127.92 19.76 128.12 19.96 ;
        RECT 127.92 15.68 128.12 15.88 ;
        RECT 127.92 11.6 128.12 11.8 ;
        RECT 128.32 56.48 128.52 56.68 ;
        RECT 128.32 52.4 128.52 52.6 ;
        RECT 128.32 48.32 128.52 48.52 ;
        RECT 128.32 44.24 128.52 44.44 ;
        RECT 128.32 40.16 128.52 40.36 ;
        RECT 128.32 36.08 128.52 36.28 ;
        RECT 128.32 32 128.52 32.2 ;
        RECT 128.32 27.92 128.52 28.12 ;
        RECT 128.32 23.84 128.52 24.04 ;
        RECT 128.32 19.76 128.52 19.96 ;
        RECT 128.32 15.68 128.52 15.88 ;
        RECT 128.32 11.6 128.52 11.8 ;
        RECT 133.44 56.48 133.64 56.68 ;
        RECT 133.44 52.4 133.64 52.6 ;
        RECT 133.44 48.32 133.64 48.52 ;
        RECT 133.44 44.24 133.64 44.44 ;
        RECT 133.44 40.16 133.64 40.36 ;
        RECT 133.44 36.08 133.64 36.28 ;
        RECT 133.44 32 133.64 32.2 ;
        RECT 133.44 27.92 133.64 28.12 ;
        RECT 133.44 23.84 133.64 24.04 ;
        RECT 133.44 19.76 133.64 19.96 ;
        RECT 133.44 15.68 133.64 15.88 ;
        RECT 133.44 11.6 133.64 11.8 ;
        RECT 133.84 56.48 134.04 56.68 ;
        RECT 133.84 52.4 134.04 52.6 ;
        RECT 133.84 48.32 134.04 48.52 ;
        RECT 133.84 44.24 134.04 44.44 ;
        RECT 133.84 40.16 134.04 40.36 ;
        RECT 133.84 36.08 134.04 36.28 ;
        RECT 133.84 32 134.04 32.2 ;
        RECT 133.84 27.92 134.04 28.12 ;
        RECT 133.84 23.84 134.04 24.04 ;
        RECT 133.84 19.76 134.04 19.96 ;
        RECT 133.84 15.68 134.04 15.88 ;
        RECT 133.84 11.6 134.04 11.8 ;
        RECT 138.96 56.48 139.16 56.68 ;
        RECT 138.96 52.4 139.16 52.6 ;
        RECT 138.96 48.32 139.16 48.52 ;
        RECT 138.96 44.24 139.16 44.44 ;
        RECT 138.96 40.16 139.16 40.36 ;
        RECT 138.96 36.08 139.16 36.28 ;
        RECT 138.96 32 139.16 32.2 ;
        RECT 138.96 27.92 139.16 28.12 ;
        RECT 138.96 23.84 139.16 24.04 ;
        RECT 138.96 19.76 139.16 19.96 ;
        RECT 138.96 15.68 139.16 15.88 ;
        RECT 138.96 11.6 139.16 11.8 ;
        RECT 139.36 56.48 139.56 56.68 ;
        RECT 139.36 52.4 139.56 52.6 ;
        RECT 139.36 48.32 139.56 48.52 ;
        RECT 139.36 44.24 139.56 44.44 ;
        RECT 139.36 40.16 139.56 40.36 ;
        RECT 139.36 36.08 139.56 36.28 ;
        RECT 139.36 32 139.56 32.2 ;
        RECT 139.36 27.92 139.56 28.12 ;
        RECT 139.36 23.84 139.56 24.04 ;
        RECT 139.36 19.76 139.56 19.96 ;
        RECT 139.36 15.68 139.56 15.88 ;
        RECT 139.36 11.6 139.56 11.8 ;
        RECT 144.48 56.48 144.68 56.68 ;
        RECT 144.48 52.4 144.68 52.6 ;
        RECT 144.48 48.32 144.68 48.52 ;
        RECT 144.48 44.24 144.68 44.44 ;
        RECT 144.48 40.16 144.68 40.36 ;
        RECT 144.48 36.08 144.68 36.28 ;
        RECT 144.48 32 144.68 32.2 ;
        RECT 144.48 27.92 144.68 28.12 ;
        RECT 144.48 23.84 144.68 24.04 ;
        RECT 144.48 19.76 144.68 19.96 ;
        RECT 144.48 15.68 144.68 15.88 ;
        RECT 144.48 11.6 144.68 11.8 ;
        RECT 144.88 56.48 145.08 56.68 ;
        RECT 144.88 52.4 145.08 52.6 ;
        RECT 144.88 48.32 145.08 48.52 ;
        RECT 144.88 44.24 145.08 44.44 ;
        RECT 144.88 40.16 145.08 40.36 ;
        RECT 144.88 36.08 145.08 36.28 ;
        RECT 144.88 32 145.08 32.2 ;
        RECT 144.88 27.92 145.08 28.12 ;
        RECT 144.88 23.84 145.08 24.04 ;
        RECT 144.88 19.76 145.08 19.96 ;
        RECT 144.88 15.68 145.08 15.88 ;
        RECT 144.88 11.6 145.08 11.8 ;
        RECT 150 56.48 150.2 56.68 ;
        RECT 150 52.4 150.2 52.6 ;
        RECT 150 48.32 150.2 48.52 ;
        RECT 150 44.24 150.2 44.44 ;
        RECT 150 40.16 150.2 40.36 ;
        RECT 150 36.08 150.2 36.28 ;
        RECT 150 32 150.2 32.2 ;
        RECT 150 27.92 150.2 28.12 ;
        RECT 150 23.84 150.2 24.04 ;
        RECT 150 19.76 150.2 19.96 ;
        RECT 150 15.68 150.2 15.88 ;
        RECT 150 11.6 150.2 11.8 ;
        RECT 150.4 56.48 150.6 56.68 ;
        RECT 150.4 52.4 150.6 52.6 ;
        RECT 150.4 48.32 150.6 48.52 ;
        RECT 150.4 44.24 150.6 44.44 ;
        RECT 150.4 40.16 150.6 40.36 ;
        RECT 150.4 36.08 150.6 36.28 ;
        RECT 150.4 32 150.6 32.2 ;
        RECT 150.4 27.92 150.6 28.12 ;
        RECT 150.4 23.84 150.6 24.04 ;
        RECT 150.4 19.76 150.6 19.96 ;
        RECT 150.4 15.68 150.6 15.88 ;
        RECT 150.4 11.6 150.6 11.8 ;
        RECT 155.52 56.48 155.72 56.68 ;
        RECT 155.52 52.4 155.72 52.6 ;
        RECT 155.52 48.32 155.72 48.52 ;
        RECT 155.52 44.24 155.72 44.44 ;
        RECT 155.52 40.16 155.72 40.36 ;
        RECT 155.52 36.08 155.72 36.28 ;
        RECT 155.52 32 155.72 32.2 ;
        RECT 155.52 27.92 155.72 28.12 ;
        RECT 155.52 23.84 155.72 24.04 ;
        RECT 155.52 19.76 155.72 19.96 ;
        RECT 155.52 15.68 155.72 15.88 ;
        RECT 155.52 11.6 155.72 11.8 ;
        RECT 155.92 56.48 156.12 56.68 ;
        RECT 155.92 52.4 156.12 52.6 ;
        RECT 155.92 48.32 156.12 48.52 ;
        RECT 155.92 44.24 156.12 44.44 ;
        RECT 155.92 40.16 156.12 40.36 ;
        RECT 155.92 36.08 156.12 36.28 ;
        RECT 155.92 32 156.12 32.2 ;
        RECT 155.92 27.92 156.12 28.12 ;
        RECT 155.92 23.84 156.12 24.04 ;
        RECT 155.92 19.76 156.12 19.96 ;
        RECT 155.92 15.68 156.12 15.88 ;
        RECT 155.92 11.6 156.12 11.8 ;
        RECT 161.04 56.48 161.24 56.68 ;
        RECT 161.04 52.4 161.24 52.6 ;
        RECT 161.04 48.32 161.24 48.52 ;
        RECT 161.04 44.24 161.24 44.44 ;
        RECT 161.04 40.16 161.24 40.36 ;
        RECT 161.04 36.08 161.24 36.28 ;
        RECT 161.04 32 161.24 32.2 ;
        RECT 161.04 27.92 161.24 28.12 ;
        RECT 161.04 23.84 161.24 24.04 ;
        RECT 161.04 19.76 161.24 19.96 ;
        RECT 161.04 15.68 161.24 15.88 ;
        RECT 161.04 11.6 161.24 11.8 ;
        RECT 161.44 56.48 161.64 56.68 ;
        RECT 161.44 52.4 161.64 52.6 ;
        RECT 161.44 48.32 161.64 48.52 ;
        RECT 161.44 44.24 161.64 44.44 ;
        RECT 161.44 40.16 161.64 40.36 ;
        RECT 161.44 36.08 161.64 36.28 ;
        RECT 161.44 32 161.64 32.2 ;
        RECT 161.44 27.92 161.64 28.12 ;
        RECT 161.44 23.84 161.64 24.04 ;
        RECT 161.44 19.76 161.64 19.96 ;
        RECT 161.44 15.68 161.64 15.88 ;
        RECT 161.44 11.6 161.64 11.8 ;
        RECT 166.56 56.48 166.76 56.68 ;
        RECT 166.56 52.4 166.76 52.6 ;
        RECT 166.56 48.32 166.76 48.52 ;
        RECT 166.56 44.24 166.76 44.44 ;
        RECT 166.56 40.16 166.76 40.36 ;
        RECT 166.56 36.08 166.76 36.28 ;
        RECT 166.56 32 166.76 32.2 ;
        RECT 166.56 27.92 166.76 28.12 ;
        RECT 166.56 23.84 166.76 24.04 ;
        RECT 166.56 19.76 166.76 19.96 ;
        RECT 166.56 15.68 166.76 15.88 ;
        RECT 166.56 11.6 166.76 11.8 ;
        RECT 166.96 56.48 167.16 56.68 ;
        RECT 166.96 52.4 167.16 52.6 ;
        RECT 166.96 48.32 167.16 48.52 ;
        RECT 166.96 44.24 167.16 44.44 ;
        RECT 166.96 40.16 167.16 40.36 ;
        RECT 166.96 36.08 167.16 36.28 ;
        RECT 166.96 32 167.16 32.2 ;
        RECT 166.96 27.92 167.16 28.12 ;
        RECT 166.96 23.84 167.16 24.04 ;
        RECT 166.96 19.76 167.16 19.96 ;
        RECT 166.96 15.68 167.16 15.88 ;
        RECT 166.96 11.6 167.16 11.8 ;
        RECT 172.08 56.48 172.28 56.68 ;
        RECT 172.08 52.4 172.28 52.6 ;
        RECT 172.08 48.32 172.28 48.52 ;
        RECT 172.08 44.24 172.28 44.44 ;
        RECT 172.08 40.16 172.28 40.36 ;
        RECT 172.08 36.08 172.28 36.28 ;
        RECT 172.08 32 172.28 32.2 ;
        RECT 172.08 27.92 172.28 28.12 ;
        RECT 172.08 23.84 172.28 24.04 ;
        RECT 172.08 19.76 172.28 19.96 ;
        RECT 172.08 15.68 172.28 15.88 ;
        RECT 172.08 11.6 172.28 11.8 ;
        RECT 172.48 56.48 172.68 56.68 ;
        RECT 172.48 52.4 172.68 52.6 ;
        RECT 172.48 48.32 172.68 48.52 ;
        RECT 172.48 44.24 172.68 44.44 ;
        RECT 172.48 40.16 172.68 40.36 ;
        RECT 172.48 36.08 172.68 36.28 ;
        RECT 172.48 32 172.68 32.2 ;
        RECT 172.48 27.92 172.68 28.12 ;
        RECT 172.48 23.84 172.68 24.04 ;
        RECT 172.48 19.76 172.68 19.96 ;
        RECT 172.48 15.68 172.68 15.88 ;
        RECT 172.48 11.6 172.68 11.8 ;
        RECT 177.6 56.48 177.8 56.68 ;
        RECT 177.6 52.4 177.8 52.6 ;
        RECT 177.6 48.32 177.8 48.52 ;
        RECT 177.6 44.24 177.8 44.44 ;
        RECT 177.6 40.16 177.8 40.36 ;
        RECT 177.6 36.08 177.8 36.28 ;
        RECT 177.6 32 177.8 32.2 ;
        RECT 177.6 27.92 177.8 28.12 ;
        RECT 177.6 23.84 177.8 24.04 ;
        RECT 177.6 19.76 177.8 19.96 ;
        RECT 177.6 15.68 177.8 15.88 ;
        RECT 177.6 11.6 177.8 11.8 ;
        RECT 178 56.48 178.2 56.68 ;
        RECT 178 52.4 178.2 52.6 ;
        RECT 178 48.32 178.2 48.52 ;
        RECT 178 44.24 178.2 44.44 ;
        RECT 178 40.16 178.2 40.36 ;
        RECT 178 36.08 178.2 36.28 ;
        RECT 178 32 178.2 32.2 ;
        RECT 178 27.92 178.2 28.12 ;
        RECT 178 23.84 178.2 24.04 ;
        RECT 178 19.76 178.2 19.96 ;
        RECT 178 15.68 178.2 15.88 ;
        RECT 178 11.6 178.2 11.8 ;
        RECT 183.12 56.48 183.32 56.68 ;
        RECT 183.12 52.4 183.32 52.6 ;
        RECT 183.12 48.32 183.32 48.52 ;
        RECT 183.12 44.24 183.32 44.44 ;
        RECT 183.12 40.16 183.32 40.36 ;
        RECT 183.12 36.08 183.32 36.28 ;
        RECT 183.12 32 183.32 32.2 ;
        RECT 183.12 27.92 183.32 28.12 ;
        RECT 183.12 23.84 183.32 24.04 ;
        RECT 183.12 19.76 183.32 19.96 ;
        RECT 183.12 15.68 183.32 15.88 ;
        RECT 183.12 11.6 183.32 11.8 ;
        RECT 183.52 56.48 183.72 56.68 ;
        RECT 183.52 52.4 183.72 52.6 ;
        RECT 183.52 48.32 183.72 48.52 ;
        RECT 183.52 44.24 183.72 44.44 ;
        RECT 183.52 40.16 183.72 40.36 ;
        RECT 183.52 36.08 183.72 36.28 ;
        RECT 183.52 32 183.72 32.2 ;
        RECT 183.52 27.92 183.72 28.12 ;
        RECT 183.52 23.84 183.72 24.04 ;
        RECT 183.52 19.76 183.72 19.96 ;
        RECT 183.52 15.68 183.72 15.88 ;
        RECT 183.52 11.6 183.72 11.8 ;
        RECT 188.64 56.48 188.84 56.68 ;
        RECT 188.64 52.4 188.84 52.6 ;
        RECT 188.64 48.32 188.84 48.52 ;
        RECT 188.64 44.24 188.84 44.44 ;
        RECT 188.64 40.16 188.84 40.36 ;
        RECT 188.64 36.08 188.84 36.28 ;
        RECT 188.64 32 188.84 32.2 ;
        RECT 188.64 27.92 188.84 28.12 ;
        RECT 188.64 23.84 188.84 24.04 ;
        RECT 188.64 19.76 188.84 19.96 ;
        RECT 188.64 15.68 188.84 15.88 ;
        RECT 188.64 11.6 188.84 11.8 ;
        RECT 189.04 56.48 189.24 56.68 ;
        RECT 189.04 52.4 189.24 52.6 ;
        RECT 189.04 48.32 189.24 48.52 ;
        RECT 189.04 44.24 189.24 44.44 ;
        RECT 189.04 40.16 189.24 40.36 ;
        RECT 189.04 36.08 189.24 36.28 ;
        RECT 189.04 32 189.24 32.2 ;
        RECT 189.04 27.92 189.24 28.12 ;
        RECT 189.04 23.84 189.24 24.04 ;
        RECT 189.04 19.76 189.24 19.96 ;
        RECT 189.04 15.68 189.24 15.88 ;
        RECT 189.04 11.6 189.24 11.8 ;
      LAYER via ;
        RECT 11.075 56.165 11.225 56.315 ;
        RECT 11.075 50.725 11.225 50.875 ;
        RECT 11.075 45.285 11.225 45.435 ;
        RECT 11.075 39.845 11.225 39.995 ;
        RECT 11.075 34.405 11.225 34.555 ;
        RECT 11.075 28.965 11.225 29.115 ;
        RECT 11.075 23.525 11.225 23.675 ;
        RECT 11.075 18.085 11.225 18.235 ;
        RECT 11.075 12.645 11.225 12.795 ;
        RECT 13.835 56.165 13.985 56.315 ;
        RECT 13.835 50.725 13.985 50.875 ;
        RECT 13.835 45.285 13.985 45.435 ;
        RECT 13.835 39.845 13.985 39.995 ;
        RECT 13.835 34.405 13.985 34.555 ;
        RECT 13.835 28.965 13.985 29.115 ;
        RECT 13.835 23.525 13.985 23.675 ;
        RECT 13.835 18.085 13.985 18.235 ;
        RECT 13.835 12.645 13.985 12.795 ;
        RECT 16.595 56.165 16.745 56.315 ;
        RECT 16.595 50.725 16.745 50.875 ;
        RECT 16.595 45.285 16.745 45.435 ;
        RECT 16.595 39.845 16.745 39.995 ;
        RECT 16.595 34.405 16.745 34.555 ;
        RECT 16.595 28.965 16.745 29.115 ;
        RECT 16.595 23.525 16.745 23.675 ;
        RECT 16.595 18.085 16.745 18.235 ;
        RECT 16.595 12.645 16.745 12.795 ;
        RECT 19.355 56.165 19.505 56.315 ;
        RECT 19.355 50.725 19.505 50.875 ;
        RECT 19.355 45.285 19.505 45.435 ;
        RECT 19.355 39.845 19.505 39.995 ;
        RECT 19.355 34.405 19.505 34.555 ;
        RECT 19.355 28.965 19.505 29.115 ;
        RECT 19.355 23.525 19.505 23.675 ;
        RECT 19.355 18.085 19.505 18.235 ;
        RECT 19.355 12.645 19.505 12.795 ;
        RECT 22.115 56.165 22.265 56.315 ;
        RECT 22.115 50.725 22.265 50.875 ;
        RECT 22.115 45.285 22.265 45.435 ;
        RECT 22.115 39.845 22.265 39.995 ;
        RECT 22.115 34.405 22.265 34.555 ;
        RECT 22.115 28.965 22.265 29.115 ;
        RECT 22.115 23.525 22.265 23.675 ;
        RECT 22.115 18.085 22.265 18.235 ;
        RECT 22.115 12.645 22.265 12.795 ;
        RECT 24.875 56.165 25.025 56.315 ;
        RECT 24.875 50.725 25.025 50.875 ;
        RECT 24.875 45.285 25.025 45.435 ;
        RECT 24.875 39.845 25.025 39.995 ;
        RECT 24.875 34.405 25.025 34.555 ;
        RECT 24.875 28.965 25.025 29.115 ;
        RECT 24.875 23.525 25.025 23.675 ;
        RECT 24.875 18.085 25.025 18.235 ;
        RECT 24.875 12.645 25.025 12.795 ;
        RECT 27.635 56.165 27.785 56.315 ;
        RECT 27.635 50.725 27.785 50.875 ;
        RECT 27.635 45.285 27.785 45.435 ;
        RECT 27.635 39.845 27.785 39.995 ;
        RECT 27.635 34.405 27.785 34.555 ;
        RECT 27.635 28.965 27.785 29.115 ;
        RECT 27.635 23.525 27.785 23.675 ;
        RECT 27.635 18.085 27.785 18.235 ;
        RECT 27.635 12.645 27.785 12.795 ;
        RECT 30.395 56.165 30.545 56.315 ;
        RECT 30.395 50.725 30.545 50.875 ;
        RECT 30.395 45.285 30.545 45.435 ;
        RECT 30.395 39.845 30.545 39.995 ;
        RECT 30.395 34.405 30.545 34.555 ;
        RECT 30.395 28.965 30.545 29.115 ;
        RECT 30.395 23.525 30.545 23.675 ;
        RECT 30.395 18.085 30.545 18.235 ;
        RECT 30.395 12.645 30.545 12.795 ;
        RECT 33.155 56.165 33.305 56.315 ;
        RECT 33.155 50.725 33.305 50.875 ;
        RECT 33.155 45.285 33.305 45.435 ;
        RECT 33.155 39.845 33.305 39.995 ;
        RECT 33.155 34.405 33.305 34.555 ;
        RECT 33.155 28.965 33.305 29.115 ;
        RECT 33.155 23.525 33.305 23.675 ;
        RECT 33.155 18.085 33.305 18.235 ;
        RECT 33.155 12.645 33.305 12.795 ;
        RECT 35.915 56.165 36.065 56.315 ;
        RECT 35.915 50.725 36.065 50.875 ;
        RECT 35.915 45.285 36.065 45.435 ;
        RECT 35.915 39.845 36.065 39.995 ;
        RECT 35.915 34.405 36.065 34.555 ;
        RECT 35.915 28.965 36.065 29.115 ;
        RECT 35.915 23.525 36.065 23.675 ;
        RECT 35.915 18.085 36.065 18.235 ;
        RECT 35.915 12.645 36.065 12.795 ;
        RECT 38.675 56.165 38.825 56.315 ;
        RECT 38.675 50.725 38.825 50.875 ;
        RECT 38.675 45.285 38.825 45.435 ;
        RECT 38.675 39.845 38.825 39.995 ;
        RECT 38.675 34.405 38.825 34.555 ;
        RECT 38.675 28.965 38.825 29.115 ;
        RECT 38.675 23.525 38.825 23.675 ;
        RECT 38.675 18.085 38.825 18.235 ;
        RECT 38.675 12.645 38.825 12.795 ;
        RECT 41.435 56.165 41.585 56.315 ;
        RECT 41.435 50.725 41.585 50.875 ;
        RECT 41.435 45.285 41.585 45.435 ;
        RECT 41.435 39.845 41.585 39.995 ;
        RECT 41.435 34.405 41.585 34.555 ;
        RECT 41.435 28.965 41.585 29.115 ;
        RECT 41.435 23.525 41.585 23.675 ;
        RECT 41.435 18.085 41.585 18.235 ;
        RECT 41.435 12.645 41.585 12.795 ;
        RECT 44.195 56.165 44.345 56.315 ;
        RECT 44.195 50.725 44.345 50.875 ;
        RECT 44.195 45.285 44.345 45.435 ;
        RECT 44.195 39.845 44.345 39.995 ;
        RECT 44.195 34.405 44.345 34.555 ;
        RECT 44.195 28.965 44.345 29.115 ;
        RECT 44.195 23.525 44.345 23.675 ;
        RECT 44.195 18.085 44.345 18.235 ;
        RECT 44.195 12.645 44.345 12.795 ;
        RECT 46.955 56.165 47.105 56.315 ;
        RECT 46.955 50.725 47.105 50.875 ;
        RECT 46.955 45.285 47.105 45.435 ;
        RECT 46.955 39.845 47.105 39.995 ;
        RECT 46.955 34.405 47.105 34.555 ;
        RECT 46.955 28.965 47.105 29.115 ;
        RECT 46.955 23.525 47.105 23.675 ;
        RECT 46.955 18.085 47.105 18.235 ;
        RECT 46.955 12.645 47.105 12.795 ;
        RECT 49.715 56.165 49.865 56.315 ;
        RECT 49.715 50.725 49.865 50.875 ;
        RECT 49.715 45.285 49.865 45.435 ;
        RECT 49.715 39.845 49.865 39.995 ;
        RECT 49.715 34.405 49.865 34.555 ;
        RECT 49.715 28.965 49.865 29.115 ;
        RECT 49.715 23.525 49.865 23.675 ;
        RECT 49.715 18.085 49.865 18.235 ;
        RECT 49.715 12.645 49.865 12.795 ;
        RECT 52.475 56.165 52.625 56.315 ;
        RECT 52.475 50.725 52.625 50.875 ;
        RECT 52.475 45.285 52.625 45.435 ;
        RECT 52.475 39.845 52.625 39.995 ;
        RECT 52.475 34.405 52.625 34.555 ;
        RECT 52.475 28.965 52.625 29.115 ;
        RECT 52.475 23.525 52.625 23.675 ;
        RECT 52.475 18.085 52.625 18.235 ;
        RECT 52.475 12.645 52.625 12.795 ;
        RECT 55.235 56.165 55.385 56.315 ;
        RECT 55.235 50.725 55.385 50.875 ;
        RECT 55.235 45.285 55.385 45.435 ;
        RECT 55.235 39.845 55.385 39.995 ;
        RECT 55.235 34.405 55.385 34.555 ;
        RECT 55.235 28.965 55.385 29.115 ;
        RECT 55.235 23.525 55.385 23.675 ;
        RECT 55.235 18.085 55.385 18.235 ;
        RECT 55.235 12.645 55.385 12.795 ;
        RECT 57.995 56.165 58.145 56.315 ;
        RECT 57.995 50.725 58.145 50.875 ;
        RECT 57.995 45.285 58.145 45.435 ;
        RECT 57.995 39.845 58.145 39.995 ;
        RECT 57.995 34.405 58.145 34.555 ;
        RECT 57.995 28.965 58.145 29.115 ;
        RECT 57.995 23.525 58.145 23.675 ;
        RECT 57.995 18.085 58.145 18.235 ;
        RECT 57.995 12.645 58.145 12.795 ;
        RECT 60.755 56.165 60.905 56.315 ;
        RECT 60.755 50.725 60.905 50.875 ;
        RECT 60.755 45.285 60.905 45.435 ;
        RECT 60.755 39.845 60.905 39.995 ;
        RECT 60.755 34.405 60.905 34.555 ;
        RECT 60.755 28.965 60.905 29.115 ;
        RECT 60.755 23.525 60.905 23.675 ;
        RECT 60.755 18.085 60.905 18.235 ;
        RECT 60.755 12.645 60.905 12.795 ;
        RECT 63.515 56.165 63.665 56.315 ;
        RECT 63.515 50.725 63.665 50.875 ;
        RECT 63.515 45.285 63.665 45.435 ;
        RECT 63.515 39.845 63.665 39.995 ;
        RECT 63.515 34.405 63.665 34.555 ;
        RECT 63.515 28.965 63.665 29.115 ;
        RECT 63.515 23.525 63.665 23.675 ;
        RECT 63.515 18.085 63.665 18.235 ;
        RECT 63.515 12.645 63.665 12.795 ;
        RECT 66.275 56.165 66.425 56.315 ;
        RECT 66.275 50.725 66.425 50.875 ;
        RECT 66.275 45.285 66.425 45.435 ;
        RECT 66.275 39.845 66.425 39.995 ;
        RECT 66.275 34.405 66.425 34.555 ;
        RECT 66.275 28.965 66.425 29.115 ;
        RECT 66.275 23.525 66.425 23.675 ;
        RECT 66.275 18.085 66.425 18.235 ;
        RECT 66.275 12.645 66.425 12.795 ;
        RECT 69.035 56.165 69.185 56.315 ;
        RECT 69.035 50.725 69.185 50.875 ;
        RECT 69.035 45.285 69.185 45.435 ;
        RECT 69.035 39.845 69.185 39.995 ;
        RECT 69.035 34.405 69.185 34.555 ;
        RECT 69.035 28.965 69.185 29.115 ;
        RECT 69.035 23.525 69.185 23.675 ;
        RECT 69.035 18.085 69.185 18.235 ;
        RECT 69.035 12.645 69.185 12.795 ;
        RECT 71.795 56.165 71.945 56.315 ;
        RECT 71.795 50.725 71.945 50.875 ;
        RECT 71.795 45.285 71.945 45.435 ;
        RECT 71.795 39.845 71.945 39.995 ;
        RECT 71.795 34.405 71.945 34.555 ;
        RECT 71.795 28.965 71.945 29.115 ;
        RECT 71.795 23.525 71.945 23.675 ;
        RECT 71.795 18.085 71.945 18.235 ;
        RECT 71.795 12.645 71.945 12.795 ;
        RECT 74.555 56.165 74.705 56.315 ;
        RECT 74.555 50.725 74.705 50.875 ;
        RECT 74.555 45.285 74.705 45.435 ;
        RECT 74.555 39.845 74.705 39.995 ;
        RECT 74.555 34.405 74.705 34.555 ;
        RECT 74.555 28.965 74.705 29.115 ;
        RECT 74.555 23.525 74.705 23.675 ;
        RECT 74.555 18.085 74.705 18.235 ;
        RECT 74.555 12.645 74.705 12.795 ;
        RECT 77.315 56.165 77.465 56.315 ;
        RECT 77.315 50.725 77.465 50.875 ;
        RECT 77.315 45.285 77.465 45.435 ;
        RECT 77.315 39.845 77.465 39.995 ;
        RECT 77.315 34.405 77.465 34.555 ;
        RECT 77.315 28.965 77.465 29.115 ;
        RECT 77.315 23.525 77.465 23.675 ;
        RECT 77.315 18.085 77.465 18.235 ;
        RECT 77.315 12.645 77.465 12.795 ;
        RECT 80.075 56.165 80.225 56.315 ;
        RECT 80.075 50.725 80.225 50.875 ;
        RECT 80.075 45.285 80.225 45.435 ;
        RECT 80.075 39.845 80.225 39.995 ;
        RECT 80.075 34.405 80.225 34.555 ;
        RECT 80.075 28.965 80.225 29.115 ;
        RECT 80.075 23.525 80.225 23.675 ;
        RECT 80.075 18.085 80.225 18.235 ;
        RECT 80.075 12.645 80.225 12.795 ;
        RECT 82.835 56.165 82.985 56.315 ;
        RECT 82.835 50.725 82.985 50.875 ;
        RECT 82.835 45.285 82.985 45.435 ;
        RECT 82.835 39.845 82.985 39.995 ;
        RECT 82.835 34.405 82.985 34.555 ;
        RECT 82.835 28.965 82.985 29.115 ;
        RECT 82.835 23.525 82.985 23.675 ;
        RECT 82.835 18.085 82.985 18.235 ;
        RECT 82.835 12.645 82.985 12.795 ;
        RECT 85.595 56.165 85.745 56.315 ;
        RECT 85.595 50.725 85.745 50.875 ;
        RECT 85.595 45.285 85.745 45.435 ;
        RECT 85.595 39.845 85.745 39.995 ;
        RECT 85.595 34.405 85.745 34.555 ;
        RECT 85.595 28.965 85.745 29.115 ;
        RECT 85.595 23.525 85.745 23.675 ;
        RECT 85.595 18.085 85.745 18.235 ;
        RECT 85.595 12.645 85.745 12.795 ;
        RECT 88.355 56.165 88.505 56.315 ;
        RECT 88.355 50.725 88.505 50.875 ;
        RECT 88.355 45.285 88.505 45.435 ;
        RECT 88.355 39.845 88.505 39.995 ;
        RECT 88.355 34.405 88.505 34.555 ;
        RECT 88.355 28.965 88.505 29.115 ;
        RECT 88.355 23.525 88.505 23.675 ;
        RECT 88.355 18.085 88.505 18.235 ;
        RECT 88.355 12.645 88.505 12.795 ;
        RECT 91.115 56.165 91.265 56.315 ;
        RECT 91.115 50.725 91.265 50.875 ;
        RECT 91.115 45.285 91.265 45.435 ;
        RECT 91.115 39.845 91.265 39.995 ;
        RECT 91.115 34.405 91.265 34.555 ;
        RECT 91.115 28.965 91.265 29.115 ;
        RECT 91.115 23.525 91.265 23.675 ;
        RECT 91.115 18.085 91.265 18.235 ;
        RECT 91.115 12.645 91.265 12.795 ;
        RECT 93.875 56.165 94.025 56.315 ;
        RECT 93.875 50.725 94.025 50.875 ;
        RECT 93.875 45.285 94.025 45.435 ;
        RECT 93.875 39.845 94.025 39.995 ;
        RECT 93.875 34.405 94.025 34.555 ;
        RECT 93.875 28.965 94.025 29.115 ;
        RECT 93.875 23.525 94.025 23.675 ;
        RECT 93.875 18.085 94.025 18.235 ;
        RECT 93.875 12.645 94.025 12.795 ;
        RECT 96.635 56.165 96.785 56.315 ;
        RECT 96.635 50.725 96.785 50.875 ;
        RECT 96.635 45.285 96.785 45.435 ;
        RECT 96.635 39.845 96.785 39.995 ;
        RECT 96.635 34.405 96.785 34.555 ;
        RECT 96.635 28.965 96.785 29.115 ;
        RECT 96.635 23.525 96.785 23.675 ;
        RECT 96.635 18.085 96.785 18.235 ;
        RECT 96.635 12.645 96.785 12.795 ;
        RECT 99.395 56.165 99.545 56.315 ;
        RECT 99.395 50.725 99.545 50.875 ;
        RECT 99.395 45.285 99.545 45.435 ;
        RECT 99.395 39.845 99.545 39.995 ;
        RECT 99.395 34.405 99.545 34.555 ;
        RECT 99.395 28.965 99.545 29.115 ;
        RECT 99.395 23.525 99.545 23.675 ;
        RECT 99.395 18.085 99.545 18.235 ;
        RECT 99.395 12.645 99.545 12.795 ;
        RECT 102.155 56.165 102.305 56.315 ;
        RECT 102.155 50.725 102.305 50.875 ;
        RECT 102.155 45.285 102.305 45.435 ;
        RECT 102.155 39.845 102.305 39.995 ;
        RECT 102.155 34.405 102.305 34.555 ;
        RECT 102.155 28.965 102.305 29.115 ;
        RECT 102.155 23.525 102.305 23.675 ;
        RECT 102.155 18.085 102.305 18.235 ;
        RECT 102.155 12.645 102.305 12.795 ;
        RECT 104.915 56.165 105.065 56.315 ;
        RECT 104.915 50.725 105.065 50.875 ;
        RECT 104.915 45.285 105.065 45.435 ;
        RECT 104.915 39.845 105.065 39.995 ;
        RECT 104.915 34.405 105.065 34.555 ;
        RECT 104.915 28.965 105.065 29.115 ;
        RECT 104.915 23.525 105.065 23.675 ;
        RECT 104.915 18.085 105.065 18.235 ;
        RECT 104.915 12.645 105.065 12.795 ;
        RECT 107.675 56.165 107.825 56.315 ;
        RECT 107.675 50.725 107.825 50.875 ;
        RECT 107.675 45.285 107.825 45.435 ;
        RECT 107.675 39.845 107.825 39.995 ;
        RECT 107.675 34.405 107.825 34.555 ;
        RECT 107.675 28.965 107.825 29.115 ;
        RECT 107.675 23.525 107.825 23.675 ;
        RECT 107.675 18.085 107.825 18.235 ;
        RECT 107.675 12.645 107.825 12.795 ;
        RECT 110.435 56.165 110.585 56.315 ;
        RECT 110.435 50.725 110.585 50.875 ;
        RECT 110.435 45.285 110.585 45.435 ;
        RECT 110.435 39.845 110.585 39.995 ;
        RECT 110.435 34.405 110.585 34.555 ;
        RECT 110.435 28.965 110.585 29.115 ;
        RECT 110.435 23.525 110.585 23.675 ;
        RECT 110.435 18.085 110.585 18.235 ;
        RECT 110.435 12.645 110.585 12.795 ;
        RECT 113.195 56.165 113.345 56.315 ;
        RECT 113.195 50.725 113.345 50.875 ;
        RECT 113.195 45.285 113.345 45.435 ;
        RECT 113.195 39.845 113.345 39.995 ;
        RECT 113.195 34.405 113.345 34.555 ;
        RECT 113.195 28.965 113.345 29.115 ;
        RECT 113.195 23.525 113.345 23.675 ;
        RECT 113.195 18.085 113.345 18.235 ;
        RECT 113.195 12.645 113.345 12.795 ;
        RECT 115.955 56.165 116.105 56.315 ;
        RECT 115.955 50.725 116.105 50.875 ;
        RECT 115.955 45.285 116.105 45.435 ;
        RECT 115.955 39.845 116.105 39.995 ;
        RECT 115.955 34.405 116.105 34.555 ;
        RECT 115.955 28.965 116.105 29.115 ;
        RECT 115.955 23.525 116.105 23.675 ;
        RECT 115.955 18.085 116.105 18.235 ;
        RECT 115.955 12.645 116.105 12.795 ;
        RECT 118.715 56.165 118.865 56.315 ;
        RECT 118.715 50.725 118.865 50.875 ;
        RECT 118.715 45.285 118.865 45.435 ;
        RECT 118.715 39.845 118.865 39.995 ;
        RECT 118.715 34.405 118.865 34.555 ;
        RECT 118.715 28.965 118.865 29.115 ;
        RECT 118.715 23.525 118.865 23.675 ;
        RECT 118.715 18.085 118.865 18.235 ;
        RECT 118.715 12.645 118.865 12.795 ;
        RECT 121.475 56.165 121.625 56.315 ;
        RECT 121.475 50.725 121.625 50.875 ;
        RECT 121.475 45.285 121.625 45.435 ;
        RECT 121.475 39.845 121.625 39.995 ;
        RECT 121.475 34.405 121.625 34.555 ;
        RECT 121.475 28.965 121.625 29.115 ;
        RECT 121.475 23.525 121.625 23.675 ;
        RECT 121.475 18.085 121.625 18.235 ;
        RECT 121.475 12.645 121.625 12.795 ;
        RECT 124.235 56.165 124.385 56.315 ;
        RECT 124.235 50.725 124.385 50.875 ;
        RECT 124.235 45.285 124.385 45.435 ;
        RECT 124.235 39.845 124.385 39.995 ;
        RECT 124.235 34.405 124.385 34.555 ;
        RECT 124.235 28.965 124.385 29.115 ;
        RECT 124.235 23.525 124.385 23.675 ;
        RECT 124.235 18.085 124.385 18.235 ;
        RECT 124.235 12.645 124.385 12.795 ;
        RECT 126.995 56.165 127.145 56.315 ;
        RECT 126.995 50.725 127.145 50.875 ;
        RECT 126.995 45.285 127.145 45.435 ;
        RECT 126.995 39.845 127.145 39.995 ;
        RECT 126.995 34.405 127.145 34.555 ;
        RECT 126.995 28.965 127.145 29.115 ;
        RECT 126.995 23.525 127.145 23.675 ;
        RECT 126.995 18.085 127.145 18.235 ;
        RECT 126.995 12.645 127.145 12.795 ;
        RECT 129.755 56.165 129.905 56.315 ;
        RECT 129.755 50.725 129.905 50.875 ;
        RECT 129.755 45.285 129.905 45.435 ;
        RECT 129.755 39.845 129.905 39.995 ;
        RECT 129.755 34.405 129.905 34.555 ;
        RECT 129.755 28.965 129.905 29.115 ;
        RECT 129.755 23.525 129.905 23.675 ;
        RECT 129.755 18.085 129.905 18.235 ;
        RECT 129.755 12.645 129.905 12.795 ;
        RECT 132.515 56.165 132.665 56.315 ;
        RECT 132.515 50.725 132.665 50.875 ;
        RECT 132.515 45.285 132.665 45.435 ;
        RECT 132.515 39.845 132.665 39.995 ;
        RECT 132.515 34.405 132.665 34.555 ;
        RECT 132.515 28.965 132.665 29.115 ;
        RECT 132.515 23.525 132.665 23.675 ;
        RECT 132.515 18.085 132.665 18.235 ;
        RECT 132.515 12.645 132.665 12.795 ;
        RECT 135.275 56.165 135.425 56.315 ;
        RECT 135.275 50.725 135.425 50.875 ;
        RECT 135.275 45.285 135.425 45.435 ;
        RECT 135.275 39.845 135.425 39.995 ;
        RECT 135.275 34.405 135.425 34.555 ;
        RECT 135.275 28.965 135.425 29.115 ;
        RECT 135.275 23.525 135.425 23.675 ;
        RECT 135.275 18.085 135.425 18.235 ;
        RECT 135.275 12.645 135.425 12.795 ;
        RECT 138.035 56.165 138.185 56.315 ;
        RECT 138.035 50.725 138.185 50.875 ;
        RECT 138.035 45.285 138.185 45.435 ;
        RECT 138.035 39.845 138.185 39.995 ;
        RECT 138.035 34.405 138.185 34.555 ;
        RECT 138.035 28.965 138.185 29.115 ;
        RECT 138.035 23.525 138.185 23.675 ;
        RECT 138.035 18.085 138.185 18.235 ;
        RECT 138.035 12.645 138.185 12.795 ;
        RECT 140.795 56.165 140.945 56.315 ;
        RECT 140.795 50.725 140.945 50.875 ;
        RECT 140.795 45.285 140.945 45.435 ;
        RECT 140.795 39.845 140.945 39.995 ;
        RECT 140.795 34.405 140.945 34.555 ;
        RECT 140.795 28.965 140.945 29.115 ;
        RECT 140.795 23.525 140.945 23.675 ;
        RECT 140.795 18.085 140.945 18.235 ;
        RECT 140.795 12.645 140.945 12.795 ;
        RECT 143.555 56.165 143.705 56.315 ;
        RECT 143.555 50.725 143.705 50.875 ;
        RECT 143.555 45.285 143.705 45.435 ;
        RECT 143.555 39.845 143.705 39.995 ;
        RECT 143.555 34.405 143.705 34.555 ;
        RECT 143.555 28.965 143.705 29.115 ;
        RECT 143.555 23.525 143.705 23.675 ;
        RECT 143.555 18.085 143.705 18.235 ;
        RECT 143.555 12.645 143.705 12.795 ;
        RECT 146.315 56.165 146.465 56.315 ;
        RECT 146.315 50.725 146.465 50.875 ;
        RECT 146.315 45.285 146.465 45.435 ;
        RECT 146.315 39.845 146.465 39.995 ;
        RECT 146.315 34.405 146.465 34.555 ;
        RECT 146.315 28.965 146.465 29.115 ;
        RECT 146.315 23.525 146.465 23.675 ;
        RECT 146.315 18.085 146.465 18.235 ;
        RECT 146.315 12.645 146.465 12.795 ;
        RECT 149.075 56.165 149.225 56.315 ;
        RECT 149.075 50.725 149.225 50.875 ;
        RECT 149.075 45.285 149.225 45.435 ;
        RECT 149.075 39.845 149.225 39.995 ;
        RECT 149.075 34.405 149.225 34.555 ;
        RECT 149.075 28.965 149.225 29.115 ;
        RECT 149.075 23.525 149.225 23.675 ;
        RECT 149.075 18.085 149.225 18.235 ;
        RECT 149.075 12.645 149.225 12.795 ;
        RECT 151.835 56.165 151.985 56.315 ;
        RECT 151.835 50.725 151.985 50.875 ;
        RECT 151.835 45.285 151.985 45.435 ;
        RECT 151.835 39.845 151.985 39.995 ;
        RECT 151.835 34.405 151.985 34.555 ;
        RECT 151.835 28.965 151.985 29.115 ;
        RECT 151.835 23.525 151.985 23.675 ;
        RECT 151.835 18.085 151.985 18.235 ;
        RECT 151.835 12.645 151.985 12.795 ;
        RECT 154.595 56.165 154.745 56.315 ;
        RECT 154.595 50.725 154.745 50.875 ;
        RECT 154.595 45.285 154.745 45.435 ;
        RECT 154.595 39.845 154.745 39.995 ;
        RECT 154.595 34.405 154.745 34.555 ;
        RECT 154.595 28.965 154.745 29.115 ;
        RECT 154.595 23.525 154.745 23.675 ;
        RECT 154.595 18.085 154.745 18.235 ;
        RECT 154.595 12.645 154.745 12.795 ;
        RECT 157.355 56.165 157.505 56.315 ;
        RECT 157.355 50.725 157.505 50.875 ;
        RECT 157.355 45.285 157.505 45.435 ;
        RECT 157.355 39.845 157.505 39.995 ;
        RECT 157.355 34.405 157.505 34.555 ;
        RECT 157.355 28.965 157.505 29.115 ;
        RECT 157.355 23.525 157.505 23.675 ;
        RECT 157.355 18.085 157.505 18.235 ;
        RECT 157.355 12.645 157.505 12.795 ;
        RECT 160.115 56.165 160.265 56.315 ;
        RECT 160.115 50.725 160.265 50.875 ;
        RECT 160.115 45.285 160.265 45.435 ;
        RECT 160.115 39.845 160.265 39.995 ;
        RECT 160.115 34.405 160.265 34.555 ;
        RECT 160.115 28.965 160.265 29.115 ;
        RECT 160.115 23.525 160.265 23.675 ;
        RECT 160.115 18.085 160.265 18.235 ;
        RECT 160.115 12.645 160.265 12.795 ;
        RECT 162.875 56.165 163.025 56.315 ;
        RECT 162.875 50.725 163.025 50.875 ;
        RECT 162.875 45.285 163.025 45.435 ;
        RECT 162.875 39.845 163.025 39.995 ;
        RECT 162.875 34.405 163.025 34.555 ;
        RECT 162.875 28.965 163.025 29.115 ;
        RECT 162.875 23.525 163.025 23.675 ;
        RECT 162.875 18.085 163.025 18.235 ;
        RECT 162.875 12.645 163.025 12.795 ;
        RECT 165.635 56.165 165.785 56.315 ;
        RECT 165.635 50.725 165.785 50.875 ;
        RECT 165.635 45.285 165.785 45.435 ;
        RECT 165.635 39.845 165.785 39.995 ;
        RECT 165.635 34.405 165.785 34.555 ;
        RECT 165.635 28.965 165.785 29.115 ;
        RECT 165.635 23.525 165.785 23.675 ;
        RECT 165.635 18.085 165.785 18.235 ;
        RECT 165.635 12.645 165.785 12.795 ;
        RECT 168.395 56.165 168.545 56.315 ;
        RECT 168.395 50.725 168.545 50.875 ;
        RECT 168.395 45.285 168.545 45.435 ;
        RECT 168.395 39.845 168.545 39.995 ;
        RECT 168.395 34.405 168.545 34.555 ;
        RECT 168.395 28.965 168.545 29.115 ;
        RECT 168.395 23.525 168.545 23.675 ;
        RECT 168.395 18.085 168.545 18.235 ;
        RECT 168.395 12.645 168.545 12.795 ;
        RECT 171.155 56.165 171.305 56.315 ;
        RECT 171.155 50.725 171.305 50.875 ;
        RECT 171.155 45.285 171.305 45.435 ;
        RECT 171.155 39.845 171.305 39.995 ;
        RECT 171.155 34.405 171.305 34.555 ;
        RECT 171.155 28.965 171.305 29.115 ;
        RECT 171.155 23.525 171.305 23.675 ;
        RECT 171.155 18.085 171.305 18.235 ;
        RECT 171.155 12.645 171.305 12.795 ;
        RECT 173.915 56.165 174.065 56.315 ;
        RECT 173.915 50.725 174.065 50.875 ;
        RECT 173.915 45.285 174.065 45.435 ;
        RECT 173.915 39.845 174.065 39.995 ;
        RECT 173.915 34.405 174.065 34.555 ;
        RECT 173.915 28.965 174.065 29.115 ;
        RECT 173.915 23.525 174.065 23.675 ;
        RECT 173.915 18.085 174.065 18.235 ;
        RECT 173.915 12.645 174.065 12.795 ;
        RECT 176.675 56.165 176.825 56.315 ;
        RECT 176.675 50.725 176.825 50.875 ;
        RECT 176.675 45.285 176.825 45.435 ;
        RECT 176.675 39.845 176.825 39.995 ;
        RECT 176.675 34.405 176.825 34.555 ;
        RECT 176.675 28.965 176.825 29.115 ;
        RECT 176.675 23.525 176.825 23.675 ;
        RECT 176.675 18.085 176.825 18.235 ;
        RECT 176.675 12.645 176.825 12.795 ;
        RECT 179.435 56.165 179.585 56.315 ;
        RECT 179.435 50.725 179.585 50.875 ;
        RECT 179.435 45.285 179.585 45.435 ;
        RECT 179.435 39.845 179.585 39.995 ;
        RECT 179.435 34.405 179.585 34.555 ;
        RECT 179.435 28.965 179.585 29.115 ;
        RECT 179.435 23.525 179.585 23.675 ;
        RECT 179.435 18.085 179.585 18.235 ;
        RECT 179.435 12.645 179.585 12.795 ;
        RECT 182.195 56.165 182.345 56.315 ;
        RECT 182.195 50.725 182.345 50.875 ;
        RECT 182.195 45.285 182.345 45.435 ;
        RECT 182.195 39.845 182.345 39.995 ;
        RECT 182.195 34.405 182.345 34.555 ;
        RECT 182.195 28.965 182.345 29.115 ;
        RECT 182.195 23.525 182.345 23.675 ;
        RECT 182.195 18.085 182.345 18.235 ;
        RECT 182.195 12.645 182.345 12.795 ;
        RECT 184.955 56.165 185.105 56.315 ;
        RECT 184.955 50.725 185.105 50.875 ;
        RECT 184.955 45.285 185.105 45.435 ;
        RECT 184.955 39.845 185.105 39.995 ;
        RECT 184.955 34.405 185.105 34.555 ;
        RECT 184.955 28.965 185.105 29.115 ;
        RECT 184.955 23.525 185.105 23.675 ;
        RECT 184.955 18.085 185.105 18.235 ;
        RECT 184.955 12.645 185.105 12.795 ;
        RECT 187.715 56.165 187.865 56.315 ;
        RECT 187.715 50.725 187.865 50.875 ;
        RECT 187.715 45.285 187.865 45.435 ;
        RECT 187.715 39.845 187.865 39.995 ;
        RECT 187.715 34.405 187.865 34.555 ;
        RECT 187.715 28.965 187.865 29.115 ;
        RECT 187.715 23.525 187.865 23.675 ;
        RECT 187.715 18.085 187.865 18.235 ;
        RECT 187.715 12.645 187.865 12.795 ;
      LAYER via4 ;
        RECT 11.9 38.5 12.7 39.3 ;
        RECT 11.9 18.1 12.7 18.9 ;
        RECT 17.42 38.5 18.22 39.3 ;
        RECT 17.42 18.1 18.22 18.9 ;
        RECT 22.94 38.5 23.74 39.3 ;
        RECT 22.94 18.1 23.74 18.9 ;
        RECT 28.46 38.5 29.26 39.3 ;
        RECT 28.46 18.1 29.26 18.9 ;
        RECT 33.98 38.5 34.78 39.3 ;
        RECT 33.98 18.1 34.78 18.9 ;
        RECT 39.5 38.5 40.3 39.3 ;
        RECT 39.5 18.1 40.3 18.9 ;
        RECT 45.02 38.5 45.82 39.3 ;
        RECT 45.02 18.1 45.82 18.9 ;
        RECT 50.54 38.5 51.34 39.3 ;
        RECT 50.54 18.1 51.34 18.9 ;
        RECT 56.06 38.5 56.86 39.3 ;
        RECT 56.06 18.1 56.86 18.9 ;
        RECT 61.58 38.5 62.38 39.3 ;
        RECT 61.58 18.1 62.38 18.9 ;
        RECT 67.1 38.5 67.9 39.3 ;
        RECT 67.1 18.1 67.9 18.9 ;
        RECT 72.62 38.5 73.42 39.3 ;
        RECT 72.62 18.1 73.42 18.9 ;
        RECT 78.14 38.5 78.94 39.3 ;
        RECT 78.14 18.1 78.94 18.9 ;
        RECT 83.66 38.5 84.46 39.3 ;
        RECT 83.66 18.1 84.46 18.9 ;
        RECT 89.18 38.5 89.98 39.3 ;
        RECT 89.18 18.1 89.98 18.9 ;
        RECT 94.7 38.5 95.5 39.3 ;
        RECT 94.7 18.1 95.5 18.9 ;
        RECT 100.22 38.5 101.02 39.3 ;
        RECT 100.22 18.1 101.02 18.9 ;
        RECT 105.74 38.5 106.54 39.3 ;
        RECT 105.74 18.1 106.54 18.9 ;
        RECT 111.26 38.5 112.06 39.3 ;
        RECT 111.26 18.1 112.06 18.9 ;
        RECT 116.78 38.5 117.58 39.3 ;
        RECT 116.78 18.1 117.58 18.9 ;
        RECT 122.3 38.5 123.1 39.3 ;
        RECT 122.3 18.1 123.1 18.9 ;
        RECT 127.82 38.5 128.62 39.3 ;
        RECT 127.82 18.1 128.62 18.9 ;
        RECT 133.34 38.5 134.14 39.3 ;
        RECT 133.34 18.1 134.14 18.9 ;
        RECT 138.86 38.5 139.66 39.3 ;
        RECT 138.86 18.1 139.66 18.9 ;
        RECT 144.38 38.5 145.18 39.3 ;
        RECT 144.38 18.1 145.18 18.9 ;
        RECT 149.9 38.5 150.7 39.3 ;
        RECT 149.9 18.1 150.7 18.9 ;
        RECT 155.42 38.5 156.22 39.3 ;
        RECT 155.42 18.1 156.22 18.9 ;
        RECT 160.94 38.5 161.74 39.3 ;
        RECT 160.94 18.1 161.74 18.9 ;
        RECT 166.46 38.5 167.26 39.3 ;
        RECT 166.46 18.1 167.26 18.9 ;
        RECT 171.98 38.5 172.78 39.3 ;
        RECT 171.98 18.1 172.78 18.9 ;
        RECT 177.5 38.5 178.3 39.3 ;
        RECT 177.5 18.1 178.3 18.9 ;
        RECT 183.02 38.5 183.82 39.3 ;
        RECT 183.02 18.1 183.82 18.9 ;
        RECT 188.54 38.5 189.34 39.3 ;
        RECT 188.54 18.1 189.34 18.9 ;
      LAYER mcon ;
        RECT 163.325 39.835 163.495 40.005 ;
        RECT 163.325 34.395 163.495 34.565 ;
        RECT 163.325 28.955 163.495 29.125 ;
        RECT 163.325 23.515 163.495 23.685 ;
        RECT 163.325 18.075 163.495 18.245 ;
        RECT 163.325 12.635 163.495 12.805 ;
        RECT 163.785 56.155 163.955 56.325 ;
        RECT 163.785 50.715 163.955 50.885 ;
        RECT 163.785 45.275 163.955 45.445 ;
        RECT 163.785 39.835 163.955 40.005 ;
        RECT 163.785 34.395 163.955 34.565 ;
        RECT 163.785 28.955 163.955 29.125 ;
        RECT 163.785 23.515 163.955 23.685 ;
        RECT 163.785 18.075 163.955 18.245 ;
        RECT 163.785 12.635 163.955 12.805 ;
        RECT 164.245 56.155 164.415 56.325 ;
        RECT 164.245 50.715 164.415 50.885 ;
        RECT 164.245 45.275 164.415 45.445 ;
        RECT 164.245 39.835 164.415 40.005 ;
        RECT 164.245 34.395 164.415 34.565 ;
        RECT 164.245 28.955 164.415 29.125 ;
        RECT 164.245 23.515 164.415 23.685 ;
        RECT 164.245 18.075 164.415 18.245 ;
        RECT 164.245 12.635 164.415 12.805 ;
        RECT 164.705 56.155 164.875 56.325 ;
        RECT 164.705 50.715 164.875 50.885 ;
        RECT 164.705 45.275 164.875 45.445 ;
        RECT 164.705 39.835 164.875 40.005 ;
        RECT 164.705 34.395 164.875 34.565 ;
        RECT 164.705 28.955 164.875 29.125 ;
        RECT 164.705 23.515 164.875 23.685 ;
        RECT 164.705 18.075 164.875 18.245 ;
        RECT 164.705 12.635 164.875 12.805 ;
        RECT 165.165 56.155 165.335 56.325 ;
        RECT 165.165 50.715 165.335 50.885 ;
        RECT 165.165 45.275 165.335 45.445 ;
        RECT 165.165 39.835 165.335 40.005 ;
        RECT 165.165 34.395 165.335 34.565 ;
        RECT 165.165 28.955 165.335 29.125 ;
        RECT 165.165 23.515 165.335 23.685 ;
        RECT 165.165 18.075 165.335 18.245 ;
        RECT 165.165 12.635 165.335 12.805 ;
        RECT 165.625 56.155 165.795 56.325 ;
        RECT 165.625 50.715 165.795 50.885 ;
        RECT 165.625 45.275 165.795 45.445 ;
        RECT 165.625 39.835 165.795 40.005 ;
        RECT 165.625 34.395 165.795 34.565 ;
        RECT 165.625 28.955 165.795 29.125 ;
        RECT 165.625 23.515 165.795 23.685 ;
        RECT 165.625 18.075 165.795 18.245 ;
        RECT 165.625 12.635 165.795 12.805 ;
        RECT 166.085 56.155 166.255 56.325 ;
        RECT 166.085 50.715 166.255 50.885 ;
        RECT 166.085 45.275 166.255 45.445 ;
        RECT 166.085 39.835 166.255 40.005 ;
        RECT 166.085 34.395 166.255 34.565 ;
        RECT 166.085 28.955 166.255 29.125 ;
        RECT 166.085 23.515 166.255 23.685 ;
        RECT 166.085 18.075 166.255 18.245 ;
        RECT 166.085 12.635 166.255 12.805 ;
        RECT 166.545 56.155 166.715 56.325 ;
        RECT 166.545 50.715 166.715 50.885 ;
        RECT 166.545 45.275 166.715 45.445 ;
        RECT 166.545 39.835 166.715 40.005 ;
        RECT 166.545 34.395 166.715 34.565 ;
        RECT 166.545 28.955 166.715 29.125 ;
        RECT 166.545 23.515 166.715 23.685 ;
        RECT 166.545 18.075 166.715 18.245 ;
        RECT 166.545 12.635 166.715 12.805 ;
        RECT 167.005 56.155 167.175 56.325 ;
        RECT 167.005 50.715 167.175 50.885 ;
        RECT 167.005 45.275 167.175 45.445 ;
        RECT 167.005 39.835 167.175 40.005 ;
        RECT 167.005 34.395 167.175 34.565 ;
        RECT 167.005 28.955 167.175 29.125 ;
        RECT 167.005 23.515 167.175 23.685 ;
        RECT 167.005 18.075 167.175 18.245 ;
        RECT 167.005 12.635 167.175 12.805 ;
        RECT 167.465 56.155 167.635 56.325 ;
        RECT 167.465 50.715 167.635 50.885 ;
        RECT 167.465 45.275 167.635 45.445 ;
        RECT 167.465 39.835 167.635 40.005 ;
        RECT 167.465 34.395 167.635 34.565 ;
        RECT 167.465 28.955 167.635 29.125 ;
        RECT 167.465 23.515 167.635 23.685 ;
        RECT 167.465 18.075 167.635 18.245 ;
        RECT 167.465 12.635 167.635 12.805 ;
        RECT 167.925 56.155 168.095 56.325 ;
        RECT 167.925 50.715 168.095 50.885 ;
        RECT 167.925 45.275 168.095 45.445 ;
        RECT 167.925 39.835 168.095 40.005 ;
        RECT 167.925 34.395 168.095 34.565 ;
        RECT 167.925 28.955 168.095 29.125 ;
        RECT 167.925 23.515 168.095 23.685 ;
        RECT 167.925 18.075 168.095 18.245 ;
        RECT 167.925 12.635 168.095 12.805 ;
        RECT 168.385 56.155 168.555 56.325 ;
        RECT 168.385 50.715 168.555 50.885 ;
        RECT 168.385 45.275 168.555 45.445 ;
        RECT 168.385 39.835 168.555 40.005 ;
        RECT 168.385 34.395 168.555 34.565 ;
        RECT 168.385 28.955 168.555 29.125 ;
        RECT 168.385 23.515 168.555 23.685 ;
        RECT 168.385 18.075 168.555 18.245 ;
        RECT 168.385 12.635 168.555 12.805 ;
        RECT 168.845 56.155 169.015 56.325 ;
        RECT 168.845 50.715 169.015 50.885 ;
        RECT 168.845 45.275 169.015 45.445 ;
        RECT 168.845 39.835 169.015 40.005 ;
        RECT 168.845 34.395 169.015 34.565 ;
        RECT 168.845 28.955 169.015 29.125 ;
        RECT 168.845 23.515 169.015 23.685 ;
        RECT 168.845 18.075 169.015 18.245 ;
        RECT 168.845 12.635 169.015 12.805 ;
        RECT 169.305 56.155 169.475 56.325 ;
        RECT 169.305 50.715 169.475 50.885 ;
        RECT 169.305 45.275 169.475 45.445 ;
        RECT 169.305 39.835 169.475 40.005 ;
        RECT 169.305 34.395 169.475 34.565 ;
        RECT 169.305 28.955 169.475 29.125 ;
        RECT 169.305 23.515 169.475 23.685 ;
        RECT 169.305 18.075 169.475 18.245 ;
        RECT 169.305 12.635 169.475 12.805 ;
        RECT 169.765 56.155 169.935 56.325 ;
        RECT 169.765 50.715 169.935 50.885 ;
        RECT 169.765 45.275 169.935 45.445 ;
        RECT 169.765 39.835 169.935 40.005 ;
        RECT 169.765 34.395 169.935 34.565 ;
        RECT 169.765 28.955 169.935 29.125 ;
        RECT 169.765 23.515 169.935 23.685 ;
        RECT 169.765 18.075 169.935 18.245 ;
        RECT 169.765 12.635 169.935 12.805 ;
        RECT 170.225 56.155 170.395 56.325 ;
        RECT 170.225 50.715 170.395 50.885 ;
        RECT 170.225 45.275 170.395 45.445 ;
        RECT 170.225 39.835 170.395 40.005 ;
        RECT 170.225 34.395 170.395 34.565 ;
        RECT 170.225 28.955 170.395 29.125 ;
        RECT 170.225 23.515 170.395 23.685 ;
        RECT 170.225 18.075 170.395 18.245 ;
        RECT 170.225 12.635 170.395 12.805 ;
        RECT 170.685 56.155 170.855 56.325 ;
        RECT 170.685 50.715 170.855 50.885 ;
        RECT 170.685 45.275 170.855 45.445 ;
        RECT 170.685 39.835 170.855 40.005 ;
        RECT 170.685 34.395 170.855 34.565 ;
        RECT 170.685 28.955 170.855 29.125 ;
        RECT 170.685 23.515 170.855 23.685 ;
        RECT 170.685 18.075 170.855 18.245 ;
        RECT 170.685 12.635 170.855 12.805 ;
        RECT 171.145 56.155 171.315 56.325 ;
        RECT 171.145 50.715 171.315 50.885 ;
        RECT 171.145 45.275 171.315 45.445 ;
        RECT 171.145 39.835 171.315 40.005 ;
        RECT 171.145 34.395 171.315 34.565 ;
        RECT 171.145 28.955 171.315 29.125 ;
        RECT 171.145 23.515 171.315 23.685 ;
        RECT 171.145 18.075 171.315 18.245 ;
        RECT 171.145 12.635 171.315 12.805 ;
        RECT 171.605 56.155 171.775 56.325 ;
        RECT 171.605 50.715 171.775 50.885 ;
        RECT 171.605 45.275 171.775 45.445 ;
        RECT 171.605 39.835 171.775 40.005 ;
        RECT 171.605 34.395 171.775 34.565 ;
        RECT 171.605 28.955 171.775 29.125 ;
        RECT 171.605 23.515 171.775 23.685 ;
        RECT 171.605 18.075 171.775 18.245 ;
        RECT 171.605 12.635 171.775 12.805 ;
        RECT 172.065 56.155 172.235 56.325 ;
        RECT 172.065 50.715 172.235 50.885 ;
        RECT 172.065 45.275 172.235 45.445 ;
        RECT 172.065 39.835 172.235 40.005 ;
        RECT 172.065 34.395 172.235 34.565 ;
        RECT 172.065 28.955 172.235 29.125 ;
        RECT 172.065 23.515 172.235 23.685 ;
        RECT 172.065 18.075 172.235 18.245 ;
        RECT 172.065 12.635 172.235 12.805 ;
        RECT 172.525 56.155 172.695 56.325 ;
        RECT 172.525 50.715 172.695 50.885 ;
        RECT 172.525 45.275 172.695 45.445 ;
        RECT 172.525 39.835 172.695 40.005 ;
        RECT 172.525 34.395 172.695 34.565 ;
        RECT 172.525 28.955 172.695 29.125 ;
        RECT 172.525 23.515 172.695 23.685 ;
        RECT 172.525 18.075 172.695 18.245 ;
        RECT 172.525 12.635 172.695 12.805 ;
        RECT 172.985 56.155 173.155 56.325 ;
        RECT 172.985 50.715 173.155 50.885 ;
        RECT 172.985 45.275 173.155 45.445 ;
        RECT 172.985 39.835 173.155 40.005 ;
        RECT 172.985 34.395 173.155 34.565 ;
        RECT 172.985 28.955 173.155 29.125 ;
        RECT 172.985 23.515 173.155 23.685 ;
        RECT 172.985 18.075 173.155 18.245 ;
        RECT 172.985 12.635 173.155 12.805 ;
        RECT 173.445 56.155 173.615 56.325 ;
        RECT 173.445 50.715 173.615 50.885 ;
        RECT 173.445 45.275 173.615 45.445 ;
        RECT 173.445 39.835 173.615 40.005 ;
        RECT 173.445 34.395 173.615 34.565 ;
        RECT 173.445 28.955 173.615 29.125 ;
        RECT 173.445 23.515 173.615 23.685 ;
        RECT 173.445 18.075 173.615 18.245 ;
        RECT 173.445 12.635 173.615 12.805 ;
        RECT 173.905 56.155 174.075 56.325 ;
        RECT 173.905 50.715 174.075 50.885 ;
        RECT 173.905 45.275 174.075 45.445 ;
        RECT 173.905 39.835 174.075 40.005 ;
        RECT 173.905 34.395 174.075 34.565 ;
        RECT 173.905 28.955 174.075 29.125 ;
        RECT 173.905 23.515 174.075 23.685 ;
        RECT 173.905 18.075 174.075 18.245 ;
        RECT 173.905 12.635 174.075 12.805 ;
        RECT 174.365 56.155 174.535 56.325 ;
        RECT 174.365 50.715 174.535 50.885 ;
        RECT 174.365 45.275 174.535 45.445 ;
        RECT 174.365 39.835 174.535 40.005 ;
        RECT 174.365 34.395 174.535 34.565 ;
        RECT 174.365 28.955 174.535 29.125 ;
        RECT 174.365 23.515 174.535 23.685 ;
        RECT 174.365 18.075 174.535 18.245 ;
        RECT 174.365 12.635 174.535 12.805 ;
        RECT 174.825 56.155 174.995 56.325 ;
        RECT 174.825 50.715 174.995 50.885 ;
        RECT 174.825 45.275 174.995 45.445 ;
        RECT 174.825 39.835 174.995 40.005 ;
        RECT 174.825 34.395 174.995 34.565 ;
        RECT 174.825 28.955 174.995 29.125 ;
        RECT 174.825 23.515 174.995 23.685 ;
        RECT 174.825 18.075 174.995 18.245 ;
        RECT 174.825 12.635 174.995 12.805 ;
        RECT 175.285 56.155 175.455 56.325 ;
        RECT 175.285 50.715 175.455 50.885 ;
        RECT 175.285 45.275 175.455 45.445 ;
        RECT 175.285 39.835 175.455 40.005 ;
        RECT 175.285 34.395 175.455 34.565 ;
        RECT 175.285 28.955 175.455 29.125 ;
        RECT 175.285 23.515 175.455 23.685 ;
        RECT 175.285 18.075 175.455 18.245 ;
        RECT 175.285 12.635 175.455 12.805 ;
        RECT 175.745 56.155 175.915 56.325 ;
        RECT 175.745 50.715 175.915 50.885 ;
        RECT 175.745 45.275 175.915 45.445 ;
        RECT 175.745 39.835 175.915 40.005 ;
        RECT 175.745 34.395 175.915 34.565 ;
        RECT 175.745 28.955 175.915 29.125 ;
        RECT 175.745 23.515 175.915 23.685 ;
        RECT 175.745 18.075 175.915 18.245 ;
        RECT 175.745 12.635 175.915 12.805 ;
        RECT 176.205 56.155 176.375 56.325 ;
        RECT 176.205 50.715 176.375 50.885 ;
        RECT 176.205 45.275 176.375 45.445 ;
        RECT 176.205 39.835 176.375 40.005 ;
        RECT 176.205 34.395 176.375 34.565 ;
        RECT 176.205 28.955 176.375 29.125 ;
        RECT 176.205 23.515 176.375 23.685 ;
        RECT 176.205 18.075 176.375 18.245 ;
        RECT 176.205 12.635 176.375 12.805 ;
        RECT 176.665 56.155 176.835 56.325 ;
        RECT 176.665 50.715 176.835 50.885 ;
        RECT 176.665 45.275 176.835 45.445 ;
        RECT 176.665 39.835 176.835 40.005 ;
        RECT 176.665 34.395 176.835 34.565 ;
        RECT 176.665 28.955 176.835 29.125 ;
        RECT 176.665 23.515 176.835 23.685 ;
        RECT 176.665 18.075 176.835 18.245 ;
        RECT 176.665 12.635 176.835 12.805 ;
        RECT 177.125 56.155 177.295 56.325 ;
        RECT 177.125 50.715 177.295 50.885 ;
        RECT 177.125 45.275 177.295 45.445 ;
        RECT 177.125 39.835 177.295 40.005 ;
        RECT 177.125 34.395 177.295 34.565 ;
        RECT 177.125 28.955 177.295 29.125 ;
        RECT 177.125 23.515 177.295 23.685 ;
        RECT 177.125 18.075 177.295 18.245 ;
        RECT 177.125 12.635 177.295 12.805 ;
        RECT 177.585 56.155 177.755 56.325 ;
        RECT 177.585 50.715 177.755 50.885 ;
        RECT 177.585 45.275 177.755 45.445 ;
        RECT 177.585 39.835 177.755 40.005 ;
        RECT 177.585 34.395 177.755 34.565 ;
        RECT 177.585 28.955 177.755 29.125 ;
        RECT 177.585 23.515 177.755 23.685 ;
        RECT 177.585 18.075 177.755 18.245 ;
        RECT 177.585 12.635 177.755 12.805 ;
        RECT 178.045 56.155 178.215 56.325 ;
        RECT 178.045 50.715 178.215 50.885 ;
        RECT 178.045 45.275 178.215 45.445 ;
        RECT 178.045 39.835 178.215 40.005 ;
        RECT 178.045 34.395 178.215 34.565 ;
        RECT 178.045 28.955 178.215 29.125 ;
        RECT 178.045 23.515 178.215 23.685 ;
        RECT 178.045 18.075 178.215 18.245 ;
        RECT 178.045 12.635 178.215 12.805 ;
        RECT 178.505 56.155 178.675 56.325 ;
        RECT 178.505 50.715 178.675 50.885 ;
        RECT 178.505 45.275 178.675 45.445 ;
        RECT 178.505 39.835 178.675 40.005 ;
        RECT 178.505 34.395 178.675 34.565 ;
        RECT 178.505 28.955 178.675 29.125 ;
        RECT 178.505 23.515 178.675 23.685 ;
        RECT 178.505 18.075 178.675 18.245 ;
        RECT 178.505 12.635 178.675 12.805 ;
        RECT 178.965 56.155 179.135 56.325 ;
        RECT 178.965 50.715 179.135 50.885 ;
        RECT 178.965 45.275 179.135 45.445 ;
        RECT 178.965 39.835 179.135 40.005 ;
        RECT 178.965 34.395 179.135 34.565 ;
        RECT 178.965 28.955 179.135 29.125 ;
        RECT 178.965 23.515 179.135 23.685 ;
        RECT 178.965 18.075 179.135 18.245 ;
        RECT 178.965 12.635 179.135 12.805 ;
        RECT 179.425 56.155 179.595 56.325 ;
        RECT 179.425 50.715 179.595 50.885 ;
        RECT 179.425 45.275 179.595 45.445 ;
        RECT 179.425 39.835 179.595 40.005 ;
        RECT 179.425 34.395 179.595 34.565 ;
        RECT 179.425 28.955 179.595 29.125 ;
        RECT 179.425 23.515 179.595 23.685 ;
        RECT 179.425 18.075 179.595 18.245 ;
        RECT 179.425 12.635 179.595 12.805 ;
        RECT 179.885 56.155 180.055 56.325 ;
        RECT 179.885 50.715 180.055 50.885 ;
        RECT 179.885 45.275 180.055 45.445 ;
        RECT 179.885 39.835 180.055 40.005 ;
        RECT 179.885 34.395 180.055 34.565 ;
        RECT 179.885 28.955 180.055 29.125 ;
        RECT 179.885 23.515 180.055 23.685 ;
        RECT 179.885 18.075 180.055 18.245 ;
        RECT 179.885 12.635 180.055 12.805 ;
        RECT 180.345 56.155 180.515 56.325 ;
        RECT 180.345 50.715 180.515 50.885 ;
        RECT 180.345 45.275 180.515 45.445 ;
        RECT 180.345 39.835 180.515 40.005 ;
        RECT 180.345 34.395 180.515 34.565 ;
        RECT 180.345 28.955 180.515 29.125 ;
        RECT 180.345 23.515 180.515 23.685 ;
        RECT 180.345 18.075 180.515 18.245 ;
        RECT 180.345 12.635 180.515 12.805 ;
        RECT 180.805 56.155 180.975 56.325 ;
        RECT 180.805 50.715 180.975 50.885 ;
        RECT 180.805 45.275 180.975 45.445 ;
        RECT 180.805 39.835 180.975 40.005 ;
        RECT 180.805 34.395 180.975 34.565 ;
        RECT 180.805 28.955 180.975 29.125 ;
        RECT 180.805 23.515 180.975 23.685 ;
        RECT 180.805 18.075 180.975 18.245 ;
        RECT 180.805 12.635 180.975 12.805 ;
        RECT 181.265 56.155 181.435 56.325 ;
        RECT 181.265 50.715 181.435 50.885 ;
        RECT 181.265 45.275 181.435 45.445 ;
        RECT 181.265 39.835 181.435 40.005 ;
        RECT 181.265 34.395 181.435 34.565 ;
        RECT 181.265 28.955 181.435 29.125 ;
        RECT 181.265 23.515 181.435 23.685 ;
        RECT 181.265 18.075 181.435 18.245 ;
        RECT 181.265 12.635 181.435 12.805 ;
        RECT 181.725 56.155 181.895 56.325 ;
        RECT 181.725 50.715 181.895 50.885 ;
        RECT 181.725 45.275 181.895 45.445 ;
        RECT 181.725 39.835 181.895 40.005 ;
        RECT 181.725 34.395 181.895 34.565 ;
        RECT 181.725 28.955 181.895 29.125 ;
        RECT 181.725 23.515 181.895 23.685 ;
        RECT 181.725 18.075 181.895 18.245 ;
        RECT 181.725 12.635 181.895 12.805 ;
        RECT 182.185 56.155 182.355 56.325 ;
        RECT 182.185 50.715 182.355 50.885 ;
        RECT 182.185 45.275 182.355 45.445 ;
        RECT 182.185 39.835 182.355 40.005 ;
        RECT 182.185 34.395 182.355 34.565 ;
        RECT 182.185 28.955 182.355 29.125 ;
        RECT 182.185 23.515 182.355 23.685 ;
        RECT 182.185 18.075 182.355 18.245 ;
        RECT 182.185 12.635 182.355 12.805 ;
        RECT 182.645 56.155 182.815 56.325 ;
        RECT 182.645 50.715 182.815 50.885 ;
        RECT 182.645 45.275 182.815 45.445 ;
        RECT 182.645 39.835 182.815 40.005 ;
        RECT 182.645 34.395 182.815 34.565 ;
        RECT 182.645 28.955 182.815 29.125 ;
        RECT 182.645 23.515 182.815 23.685 ;
        RECT 182.645 18.075 182.815 18.245 ;
        RECT 182.645 12.635 182.815 12.805 ;
        RECT 183.105 56.155 183.275 56.325 ;
        RECT 183.105 50.715 183.275 50.885 ;
        RECT 183.105 45.275 183.275 45.445 ;
        RECT 183.105 39.835 183.275 40.005 ;
        RECT 183.105 34.395 183.275 34.565 ;
        RECT 183.105 28.955 183.275 29.125 ;
        RECT 183.105 23.515 183.275 23.685 ;
        RECT 183.105 18.075 183.275 18.245 ;
        RECT 183.105 12.635 183.275 12.805 ;
        RECT 183.565 56.155 183.735 56.325 ;
        RECT 183.565 50.715 183.735 50.885 ;
        RECT 183.565 45.275 183.735 45.445 ;
        RECT 183.565 39.835 183.735 40.005 ;
        RECT 183.565 34.395 183.735 34.565 ;
        RECT 183.565 28.955 183.735 29.125 ;
        RECT 183.565 23.515 183.735 23.685 ;
        RECT 183.565 18.075 183.735 18.245 ;
        RECT 183.565 12.635 183.735 12.805 ;
        RECT 184.025 56.155 184.195 56.325 ;
        RECT 184.025 50.715 184.195 50.885 ;
        RECT 184.025 45.275 184.195 45.445 ;
        RECT 184.025 39.835 184.195 40.005 ;
        RECT 184.025 34.395 184.195 34.565 ;
        RECT 184.025 28.955 184.195 29.125 ;
        RECT 184.025 23.515 184.195 23.685 ;
        RECT 184.025 18.075 184.195 18.245 ;
        RECT 184.025 12.635 184.195 12.805 ;
        RECT 184.485 56.155 184.655 56.325 ;
        RECT 184.485 50.715 184.655 50.885 ;
        RECT 184.485 45.275 184.655 45.445 ;
        RECT 184.485 39.835 184.655 40.005 ;
        RECT 184.485 34.395 184.655 34.565 ;
        RECT 184.485 28.955 184.655 29.125 ;
        RECT 184.485 23.515 184.655 23.685 ;
        RECT 184.485 18.075 184.655 18.245 ;
        RECT 184.485 12.635 184.655 12.805 ;
        RECT 184.945 56.155 185.115 56.325 ;
        RECT 184.945 50.715 185.115 50.885 ;
        RECT 184.945 45.275 185.115 45.445 ;
        RECT 184.945 39.835 185.115 40.005 ;
        RECT 184.945 34.395 185.115 34.565 ;
        RECT 184.945 28.955 185.115 29.125 ;
        RECT 184.945 23.515 185.115 23.685 ;
        RECT 184.945 18.075 185.115 18.245 ;
        RECT 184.945 12.635 185.115 12.805 ;
        RECT 185.405 56.155 185.575 56.325 ;
        RECT 185.405 50.715 185.575 50.885 ;
        RECT 185.405 45.275 185.575 45.445 ;
        RECT 185.405 39.835 185.575 40.005 ;
        RECT 185.405 34.395 185.575 34.565 ;
        RECT 185.405 28.955 185.575 29.125 ;
        RECT 185.405 23.515 185.575 23.685 ;
        RECT 185.405 18.075 185.575 18.245 ;
        RECT 185.405 12.635 185.575 12.805 ;
        RECT 185.865 56.155 186.035 56.325 ;
        RECT 185.865 50.715 186.035 50.885 ;
        RECT 185.865 45.275 186.035 45.445 ;
        RECT 185.865 39.835 186.035 40.005 ;
        RECT 185.865 34.395 186.035 34.565 ;
        RECT 185.865 28.955 186.035 29.125 ;
        RECT 185.865 23.515 186.035 23.685 ;
        RECT 185.865 18.075 186.035 18.245 ;
        RECT 185.865 12.635 186.035 12.805 ;
        RECT 186.325 56.155 186.495 56.325 ;
        RECT 186.325 50.715 186.495 50.885 ;
        RECT 186.325 45.275 186.495 45.445 ;
        RECT 186.325 39.835 186.495 40.005 ;
        RECT 186.325 34.395 186.495 34.565 ;
        RECT 186.325 28.955 186.495 29.125 ;
        RECT 186.325 23.515 186.495 23.685 ;
        RECT 186.325 18.075 186.495 18.245 ;
        RECT 186.325 12.635 186.495 12.805 ;
        RECT 186.785 56.155 186.955 56.325 ;
        RECT 186.785 50.715 186.955 50.885 ;
        RECT 186.785 45.275 186.955 45.445 ;
        RECT 186.785 39.835 186.955 40.005 ;
        RECT 186.785 34.395 186.955 34.565 ;
        RECT 186.785 28.955 186.955 29.125 ;
        RECT 186.785 23.515 186.955 23.685 ;
        RECT 186.785 18.075 186.955 18.245 ;
        RECT 186.785 12.635 186.955 12.805 ;
        RECT 187.245 56.155 187.415 56.325 ;
        RECT 187.245 50.715 187.415 50.885 ;
        RECT 187.245 45.275 187.415 45.445 ;
        RECT 187.245 39.835 187.415 40.005 ;
        RECT 187.245 34.395 187.415 34.565 ;
        RECT 187.245 28.955 187.415 29.125 ;
        RECT 187.245 23.515 187.415 23.685 ;
        RECT 187.245 18.075 187.415 18.245 ;
        RECT 187.245 12.635 187.415 12.805 ;
        RECT 187.705 56.155 187.875 56.325 ;
        RECT 187.705 50.715 187.875 50.885 ;
        RECT 187.705 45.275 187.875 45.445 ;
        RECT 187.705 39.835 187.875 40.005 ;
        RECT 187.705 34.395 187.875 34.565 ;
        RECT 187.705 28.955 187.875 29.125 ;
        RECT 187.705 23.515 187.875 23.685 ;
        RECT 187.705 18.075 187.875 18.245 ;
        RECT 187.705 12.635 187.875 12.805 ;
        RECT 188.165 56.155 188.335 56.325 ;
        RECT 188.165 50.715 188.335 50.885 ;
        RECT 188.165 45.275 188.335 45.445 ;
        RECT 188.165 39.835 188.335 40.005 ;
        RECT 188.165 34.395 188.335 34.565 ;
        RECT 188.165 28.955 188.335 29.125 ;
        RECT 188.165 23.515 188.335 23.685 ;
        RECT 188.165 18.075 188.335 18.245 ;
        RECT 188.165 12.635 188.335 12.805 ;
        RECT 188.625 56.155 188.795 56.325 ;
        RECT 188.625 50.715 188.795 50.885 ;
        RECT 188.625 45.275 188.795 45.445 ;
        RECT 188.625 39.835 188.795 40.005 ;
        RECT 188.625 34.395 188.795 34.565 ;
        RECT 188.625 28.955 188.795 29.125 ;
        RECT 188.625 23.515 188.795 23.685 ;
        RECT 188.625 18.075 188.795 18.245 ;
        RECT 188.625 12.635 188.795 12.805 ;
        RECT 189.085 56.155 189.255 56.325 ;
        RECT 189.085 50.715 189.255 50.885 ;
        RECT 189.085 45.275 189.255 45.445 ;
        RECT 189.085 39.835 189.255 40.005 ;
        RECT 189.085 34.395 189.255 34.565 ;
        RECT 189.085 28.955 189.255 29.125 ;
        RECT 189.085 23.515 189.255 23.685 ;
        RECT 189.085 18.075 189.255 18.245 ;
        RECT 189.085 12.635 189.255 12.805 ;
        RECT 189.545 56.155 189.715 56.325 ;
        RECT 189.545 50.715 189.715 50.885 ;
        RECT 189.545 45.275 189.715 45.445 ;
        RECT 189.545 39.835 189.715 40.005 ;
        RECT 189.545 34.395 189.715 34.565 ;
        RECT 189.545 28.955 189.715 29.125 ;
        RECT 189.545 23.515 189.715 23.685 ;
        RECT 189.545 18.075 189.715 18.245 ;
        RECT 189.545 12.635 189.715 12.805 ;
        RECT 112.265 45.275 112.435 45.445 ;
        RECT 112.265 39.835 112.435 40.005 ;
        RECT 112.265 34.395 112.435 34.565 ;
        RECT 112.265 28.955 112.435 29.125 ;
        RECT 112.265 23.515 112.435 23.685 ;
        RECT 112.265 18.075 112.435 18.245 ;
        RECT 112.265 12.635 112.435 12.805 ;
        RECT 112.725 56.155 112.895 56.325 ;
        RECT 112.725 50.715 112.895 50.885 ;
        RECT 112.725 45.275 112.895 45.445 ;
        RECT 112.725 39.835 112.895 40.005 ;
        RECT 112.725 34.395 112.895 34.565 ;
        RECT 112.725 28.955 112.895 29.125 ;
        RECT 112.725 23.515 112.895 23.685 ;
        RECT 112.725 18.075 112.895 18.245 ;
        RECT 112.725 12.635 112.895 12.805 ;
        RECT 113.185 56.155 113.355 56.325 ;
        RECT 113.185 50.715 113.355 50.885 ;
        RECT 113.185 45.275 113.355 45.445 ;
        RECT 113.185 39.835 113.355 40.005 ;
        RECT 113.185 34.395 113.355 34.565 ;
        RECT 113.185 28.955 113.355 29.125 ;
        RECT 113.185 23.515 113.355 23.685 ;
        RECT 113.185 18.075 113.355 18.245 ;
        RECT 113.185 12.635 113.355 12.805 ;
        RECT 113.645 56.155 113.815 56.325 ;
        RECT 113.645 50.715 113.815 50.885 ;
        RECT 113.645 45.275 113.815 45.445 ;
        RECT 113.645 39.835 113.815 40.005 ;
        RECT 113.645 34.395 113.815 34.565 ;
        RECT 113.645 28.955 113.815 29.125 ;
        RECT 113.645 23.515 113.815 23.685 ;
        RECT 113.645 18.075 113.815 18.245 ;
        RECT 113.645 12.635 113.815 12.805 ;
        RECT 114.105 56.155 114.275 56.325 ;
        RECT 114.105 50.715 114.275 50.885 ;
        RECT 114.105 45.275 114.275 45.445 ;
        RECT 114.105 39.835 114.275 40.005 ;
        RECT 114.105 34.395 114.275 34.565 ;
        RECT 114.105 28.955 114.275 29.125 ;
        RECT 114.105 23.515 114.275 23.685 ;
        RECT 114.105 18.075 114.275 18.245 ;
        RECT 114.105 12.635 114.275 12.805 ;
        RECT 114.565 56.155 114.735 56.325 ;
        RECT 114.565 50.715 114.735 50.885 ;
        RECT 114.565 45.275 114.735 45.445 ;
        RECT 114.565 39.835 114.735 40.005 ;
        RECT 114.565 34.395 114.735 34.565 ;
        RECT 114.565 28.955 114.735 29.125 ;
        RECT 114.565 23.515 114.735 23.685 ;
        RECT 114.565 18.075 114.735 18.245 ;
        RECT 114.565 12.635 114.735 12.805 ;
        RECT 115.025 56.155 115.195 56.325 ;
        RECT 115.025 50.715 115.195 50.885 ;
        RECT 115.025 45.275 115.195 45.445 ;
        RECT 115.025 39.835 115.195 40.005 ;
        RECT 115.025 34.395 115.195 34.565 ;
        RECT 115.025 28.955 115.195 29.125 ;
        RECT 115.025 23.515 115.195 23.685 ;
        RECT 115.025 18.075 115.195 18.245 ;
        RECT 115.025 12.635 115.195 12.805 ;
        RECT 115.485 56.155 115.655 56.325 ;
        RECT 115.485 50.715 115.655 50.885 ;
        RECT 115.485 45.275 115.655 45.445 ;
        RECT 115.485 39.835 115.655 40.005 ;
        RECT 115.485 34.395 115.655 34.565 ;
        RECT 115.485 28.955 115.655 29.125 ;
        RECT 115.485 23.515 115.655 23.685 ;
        RECT 115.485 18.075 115.655 18.245 ;
        RECT 115.485 12.635 115.655 12.805 ;
        RECT 115.945 56.155 116.115 56.325 ;
        RECT 115.945 50.715 116.115 50.885 ;
        RECT 115.945 45.275 116.115 45.445 ;
        RECT 115.945 39.835 116.115 40.005 ;
        RECT 115.945 34.395 116.115 34.565 ;
        RECT 115.945 28.955 116.115 29.125 ;
        RECT 115.945 23.515 116.115 23.685 ;
        RECT 115.945 18.075 116.115 18.245 ;
        RECT 115.945 12.635 116.115 12.805 ;
        RECT 116.405 56.155 116.575 56.325 ;
        RECT 116.405 50.715 116.575 50.885 ;
        RECT 116.405 45.275 116.575 45.445 ;
        RECT 116.405 39.835 116.575 40.005 ;
        RECT 116.405 34.395 116.575 34.565 ;
        RECT 116.405 28.955 116.575 29.125 ;
        RECT 116.405 23.515 116.575 23.685 ;
        RECT 116.405 18.075 116.575 18.245 ;
        RECT 116.405 12.635 116.575 12.805 ;
        RECT 116.865 56.155 117.035 56.325 ;
        RECT 116.865 50.715 117.035 50.885 ;
        RECT 116.865 45.275 117.035 45.445 ;
        RECT 116.865 39.835 117.035 40.005 ;
        RECT 116.865 34.395 117.035 34.565 ;
        RECT 116.865 28.955 117.035 29.125 ;
        RECT 116.865 23.515 117.035 23.685 ;
        RECT 116.865 18.075 117.035 18.245 ;
        RECT 116.865 12.635 117.035 12.805 ;
        RECT 117.325 56.155 117.495 56.325 ;
        RECT 117.325 50.715 117.495 50.885 ;
        RECT 117.325 45.275 117.495 45.445 ;
        RECT 117.325 39.835 117.495 40.005 ;
        RECT 117.325 34.395 117.495 34.565 ;
        RECT 117.325 28.955 117.495 29.125 ;
        RECT 117.325 23.515 117.495 23.685 ;
        RECT 117.325 18.075 117.495 18.245 ;
        RECT 117.325 12.635 117.495 12.805 ;
        RECT 117.785 56.155 117.955 56.325 ;
        RECT 117.785 50.715 117.955 50.885 ;
        RECT 117.785 45.275 117.955 45.445 ;
        RECT 117.785 39.835 117.955 40.005 ;
        RECT 117.785 34.395 117.955 34.565 ;
        RECT 117.785 28.955 117.955 29.125 ;
        RECT 117.785 23.515 117.955 23.685 ;
        RECT 117.785 18.075 117.955 18.245 ;
        RECT 117.785 12.635 117.955 12.805 ;
        RECT 118.245 56.155 118.415 56.325 ;
        RECT 118.245 50.715 118.415 50.885 ;
        RECT 118.245 45.275 118.415 45.445 ;
        RECT 118.245 39.835 118.415 40.005 ;
        RECT 118.245 34.395 118.415 34.565 ;
        RECT 118.245 28.955 118.415 29.125 ;
        RECT 118.245 23.515 118.415 23.685 ;
        RECT 118.245 18.075 118.415 18.245 ;
        RECT 118.245 12.635 118.415 12.805 ;
        RECT 118.705 56.155 118.875 56.325 ;
        RECT 118.705 50.715 118.875 50.885 ;
        RECT 118.705 45.275 118.875 45.445 ;
        RECT 118.705 39.835 118.875 40.005 ;
        RECT 118.705 34.395 118.875 34.565 ;
        RECT 118.705 28.955 118.875 29.125 ;
        RECT 118.705 23.515 118.875 23.685 ;
        RECT 118.705 18.075 118.875 18.245 ;
        RECT 118.705 12.635 118.875 12.805 ;
        RECT 119.165 56.155 119.335 56.325 ;
        RECT 119.165 50.715 119.335 50.885 ;
        RECT 119.165 45.275 119.335 45.445 ;
        RECT 119.165 39.835 119.335 40.005 ;
        RECT 119.165 34.395 119.335 34.565 ;
        RECT 119.165 28.955 119.335 29.125 ;
        RECT 119.165 23.515 119.335 23.685 ;
        RECT 119.165 18.075 119.335 18.245 ;
        RECT 119.165 12.635 119.335 12.805 ;
        RECT 119.625 56.155 119.795 56.325 ;
        RECT 119.625 50.715 119.795 50.885 ;
        RECT 119.625 45.275 119.795 45.445 ;
        RECT 119.625 39.835 119.795 40.005 ;
        RECT 119.625 34.395 119.795 34.565 ;
        RECT 119.625 28.955 119.795 29.125 ;
        RECT 119.625 23.515 119.795 23.685 ;
        RECT 119.625 18.075 119.795 18.245 ;
        RECT 119.625 12.635 119.795 12.805 ;
        RECT 120.085 56.155 120.255 56.325 ;
        RECT 120.085 50.715 120.255 50.885 ;
        RECT 120.085 45.275 120.255 45.445 ;
        RECT 120.085 39.835 120.255 40.005 ;
        RECT 120.085 34.395 120.255 34.565 ;
        RECT 120.085 28.955 120.255 29.125 ;
        RECT 120.085 23.515 120.255 23.685 ;
        RECT 120.085 18.075 120.255 18.245 ;
        RECT 120.085 12.635 120.255 12.805 ;
        RECT 120.545 56.155 120.715 56.325 ;
        RECT 120.545 50.715 120.715 50.885 ;
        RECT 120.545 45.275 120.715 45.445 ;
        RECT 120.545 39.835 120.715 40.005 ;
        RECT 120.545 34.395 120.715 34.565 ;
        RECT 120.545 28.955 120.715 29.125 ;
        RECT 120.545 23.515 120.715 23.685 ;
        RECT 120.545 18.075 120.715 18.245 ;
        RECT 120.545 12.635 120.715 12.805 ;
        RECT 121.005 56.155 121.175 56.325 ;
        RECT 121.005 50.715 121.175 50.885 ;
        RECT 121.005 45.275 121.175 45.445 ;
        RECT 121.005 39.835 121.175 40.005 ;
        RECT 121.005 34.395 121.175 34.565 ;
        RECT 121.005 28.955 121.175 29.125 ;
        RECT 121.005 23.515 121.175 23.685 ;
        RECT 121.005 18.075 121.175 18.245 ;
        RECT 121.005 12.635 121.175 12.805 ;
        RECT 121.465 56.155 121.635 56.325 ;
        RECT 121.465 50.715 121.635 50.885 ;
        RECT 121.465 45.275 121.635 45.445 ;
        RECT 121.465 39.835 121.635 40.005 ;
        RECT 121.465 34.395 121.635 34.565 ;
        RECT 121.465 28.955 121.635 29.125 ;
        RECT 121.465 23.515 121.635 23.685 ;
        RECT 121.465 18.075 121.635 18.245 ;
        RECT 121.465 12.635 121.635 12.805 ;
        RECT 121.925 56.155 122.095 56.325 ;
        RECT 121.925 50.715 122.095 50.885 ;
        RECT 121.925 45.275 122.095 45.445 ;
        RECT 121.925 39.835 122.095 40.005 ;
        RECT 121.925 34.395 122.095 34.565 ;
        RECT 121.925 28.955 122.095 29.125 ;
        RECT 121.925 23.515 122.095 23.685 ;
        RECT 121.925 18.075 122.095 18.245 ;
        RECT 121.925 12.635 122.095 12.805 ;
        RECT 122.385 56.155 122.555 56.325 ;
        RECT 122.385 50.715 122.555 50.885 ;
        RECT 122.385 45.275 122.555 45.445 ;
        RECT 122.385 39.835 122.555 40.005 ;
        RECT 122.385 34.395 122.555 34.565 ;
        RECT 122.385 28.955 122.555 29.125 ;
        RECT 122.385 23.515 122.555 23.685 ;
        RECT 122.385 18.075 122.555 18.245 ;
        RECT 122.385 12.635 122.555 12.805 ;
        RECT 122.845 56.155 123.015 56.325 ;
        RECT 122.845 50.715 123.015 50.885 ;
        RECT 122.845 45.275 123.015 45.445 ;
        RECT 122.845 39.835 123.015 40.005 ;
        RECT 122.845 34.395 123.015 34.565 ;
        RECT 122.845 28.955 123.015 29.125 ;
        RECT 122.845 23.515 123.015 23.685 ;
        RECT 122.845 18.075 123.015 18.245 ;
        RECT 122.845 12.635 123.015 12.805 ;
        RECT 123.305 56.155 123.475 56.325 ;
        RECT 123.305 50.715 123.475 50.885 ;
        RECT 123.305 45.275 123.475 45.445 ;
        RECT 123.305 39.835 123.475 40.005 ;
        RECT 123.305 34.395 123.475 34.565 ;
        RECT 123.305 28.955 123.475 29.125 ;
        RECT 123.305 23.515 123.475 23.685 ;
        RECT 123.305 18.075 123.475 18.245 ;
        RECT 123.305 12.635 123.475 12.805 ;
        RECT 123.765 56.155 123.935 56.325 ;
        RECT 123.765 50.715 123.935 50.885 ;
        RECT 123.765 45.275 123.935 45.445 ;
        RECT 123.765 39.835 123.935 40.005 ;
        RECT 123.765 34.395 123.935 34.565 ;
        RECT 123.765 28.955 123.935 29.125 ;
        RECT 123.765 23.515 123.935 23.685 ;
        RECT 123.765 18.075 123.935 18.245 ;
        RECT 123.765 12.635 123.935 12.805 ;
        RECT 124.225 56.155 124.395 56.325 ;
        RECT 124.225 50.715 124.395 50.885 ;
        RECT 124.225 45.275 124.395 45.445 ;
        RECT 124.225 39.835 124.395 40.005 ;
        RECT 124.225 34.395 124.395 34.565 ;
        RECT 124.225 28.955 124.395 29.125 ;
        RECT 124.225 23.515 124.395 23.685 ;
        RECT 124.225 18.075 124.395 18.245 ;
        RECT 124.225 12.635 124.395 12.805 ;
        RECT 124.685 56.155 124.855 56.325 ;
        RECT 124.685 50.715 124.855 50.885 ;
        RECT 124.685 45.275 124.855 45.445 ;
        RECT 124.685 39.835 124.855 40.005 ;
        RECT 124.685 34.395 124.855 34.565 ;
        RECT 124.685 28.955 124.855 29.125 ;
        RECT 124.685 23.515 124.855 23.685 ;
        RECT 124.685 18.075 124.855 18.245 ;
        RECT 124.685 12.635 124.855 12.805 ;
        RECT 125.145 56.155 125.315 56.325 ;
        RECT 125.145 50.715 125.315 50.885 ;
        RECT 125.145 45.275 125.315 45.445 ;
        RECT 125.145 39.835 125.315 40.005 ;
        RECT 125.145 34.395 125.315 34.565 ;
        RECT 125.145 28.955 125.315 29.125 ;
        RECT 125.145 23.515 125.315 23.685 ;
        RECT 125.145 18.075 125.315 18.245 ;
        RECT 125.145 12.635 125.315 12.805 ;
        RECT 125.605 56.155 125.775 56.325 ;
        RECT 125.605 50.715 125.775 50.885 ;
        RECT 125.605 45.275 125.775 45.445 ;
        RECT 125.605 39.835 125.775 40.005 ;
        RECT 125.605 34.395 125.775 34.565 ;
        RECT 125.605 28.955 125.775 29.125 ;
        RECT 125.605 23.515 125.775 23.685 ;
        RECT 125.605 18.075 125.775 18.245 ;
        RECT 125.605 12.635 125.775 12.805 ;
        RECT 126.065 56.155 126.235 56.325 ;
        RECT 126.065 50.715 126.235 50.885 ;
        RECT 126.065 45.275 126.235 45.445 ;
        RECT 126.065 39.835 126.235 40.005 ;
        RECT 126.065 34.395 126.235 34.565 ;
        RECT 126.065 28.955 126.235 29.125 ;
        RECT 126.065 23.515 126.235 23.685 ;
        RECT 126.065 18.075 126.235 18.245 ;
        RECT 126.065 12.635 126.235 12.805 ;
        RECT 126.525 56.155 126.695 56.325 ;
        RECT 126.525 50.715 126.695 50.885 ;
        RECT 126.525 45.275 126.695 45.445 ;
        RECT 126.525 39.835 126.695 40.005 ;
        RECT 126.525 34.395 126.695 34.565 ;
        RECT 126.525 28.955 126.695 29.125 ;
        RECT 126.525 23.515 126.695 23.685 ;
        RECT 126.525 18.075 126.695 18.245 ;
        RECT 126.525 12.635 126.695 12.805 ;
        RECT 126.985 56.155 127.155 56.325 ;
        RECT 126.985 50.715 127.155 50.885 ;
        RECT 126.985 45.275 127.155 45.445 ;
        RECT 126.985 39.835 127.155 40.005 ;
        RECT 126.985 34.395 127.155 34.565 ;
        RECT 126.985 28.955 127.155 29.125 ;
        RECT 126.985 23.515 127.155 23.685 ;
        RECT 126.985 18.075 127.155 18.245 ;
        RECT 126.985 12.635 127.155 12.805 ;
        RECT 127.445 56.155 127.615 56.325 ;
        RECT 127.445 50.715 127.615 50.885 ;
        RECT 127.445 45.275 127.615 45.445 ;
        RECT 127.445 39.835 127.615 40.005 ;
        RECT 127.445 34.395 127.615 34.565 ;
        RECT 127.445 28.955 127.615 29.125 ;
        RECT 127.445 23.515 127.615 23.685 ;
        RECT 127.445 18.075 127.615 18.245 ;
        RECT 127.445 12.635 127.615 12.805 ;
        RECT 127.905 56.155 128.075 56.325 ;
        RECT 127.905 50.715 128.075 50.885 ;
        RECT 127.905 45.275 128.075 45.445 ;
        RECT 127.905 39.835 128.075 40.005 ;
        RECT 127.905 34.395 128.075 34.565 ;
        RECT 127.905 28.955 128.075 29.125 ;
        RECT 127.905 23.515 128.075 23.685 ;
        RECT 127.905 18.075 128.075 18.245 ;
        RECT 127.905 12.635 128.075 12.805 ;
        RECT 128.365 56.155 128.535 56.325 ;
        RECT 128.365 50.715 128.535 50.885 ;
        RECT 128.365 45.275 128.535 45.445 ;
        RECT 128.365 39.835 128.535 40.005 ;
        RECT 128.365 34.395 128.535 34.565 ;
        RECT 128.365 28.955 128.535 29.125 ;
        RECT 128.365 23.515 128.535 23.685 ;
        RECT 128.365 18.075 128.535 18.245 ;
        RECT 128.365 12.635 128.535 12.805 ;
        RECT 128.825 56.155 128.995 56.325 ;
        RECT 128.825 50.715 128.995 50.885 ;
        RECT 128.825 45.275 128.995 45.445 ;
        RECT 128.825 39.835 128.995 40.005 ;
        RECT 128.825 34.395 128.995 34.565 ;
        RECT 128.825 28.955 128.995 29.125 ;
        RECT 128.825 23.515 128.995 23.685 ;
        RECT 128.825 18.075 128.995 18.245 ;
        RECT 128.825 12.635 128.995 12.805 ;
        RECT 129.285 56.155 129.455 56.325 ;
        RECT 129.285 50.715 129.455 50.885 ;
        RECT 129.285 45.275 129.455 45.445 ;
        RECT 129.285 39.835 129.455 40.005 ;
        RECT 129.285 34.395 129.455 34.565 ;
        RECT 129.285 28.955 129.455 29.125 ;
        RECT 129.285 23.515 129.455 23.685 ;
        RECT 129.285 18.075 129.455 18.245 ;
        RECT 129.285 12.635 129.455 12.805 ;
        RECT 129.745 56.155 129.915 56.325 ;
        RECT 129.745 50.715 129.915 50.885 ;
        RECT 129.745 45.275 129.915 45.445 ;
        RECT 129.745 39.835 129.915 40.005 ;
        RECT 129.745 34.395 129.915 34.565 ;
        RECT 129.745 28.955 129.915 29.125 ;
        RECT 129.745 23.515 129.915 23.685 ;
        RECT 129.745 18.075 129.915 18.245 ;
        RECT 129.745 12.635 129.915 12.805 ;
        RECT 130.205 56.155 130.375 56.325 ;
        RECT 130.205 50.715 130.375 50.885 ;
        RECT 130.205 45.275 130.375 45.445 ;
        RECT 130.205 39.835 130.375 40.005 ;
        RECT 130.205 34.395 130.375 34.565 ;
        RECT 130.205 28.955 130.375 29.125 ;
        RECT 130.205 23.515 130.375 23.685 ;
        RECT 130.205 18.075 130.375 18.245 ;
        RECT 130.205 12.635 130.375 12.805 ;
        RECT 130.665 56.155 130.835 56.325 ;
        RECT 130.665 50.715 130.835 50.885 ;
        RECT 130.665 45.275 130.835 45.445 ;
        RECT 130.665 39.835 130.835 40.005 ;
        RECT 130.665 34.395 130.835 34.565 ;
        RECT 130.665 28.955 130.835 29.125 ;
        RECT 130.665 23.515 130.835 23.685 ;
        RECT 130.665 18.075 130.835 18.245 ;
        RECT 130.665 12.635 130.835 12.805 ;
        RECT 131.125 56.155 131.295 56.325 ;
        RECT 131.125 50.715 131.295 50.885 ;
        RECT 131.125 45.275 131.295 45.445 ;
        RECT 131.125 39.835 131.295 40.005 ;
        RECT 131.125 34.395 131.295 34.565 ;
        RECT 131.125 28.955 131.295 29.125 ;
        RECT 131.125 23.515 131.295 23.685 ;
        RECT 131.125 18.075 131.295 18.245 ;
        RECT 131.125 12.635 131.295 12.805 ;
        RECT 131.585 56.155 131.755 56.325 ;
        RECT 131.585 50.715 131.755 50.885 ;
        RECT 131.585 45.275 131.755 45.445 ;
        RECT 131.585 39.835 131.755 40.005 ;
        RECT 131.585 34.395 131.755 34.565 ;
        RECT 131.585 28.955 131.755 29.125 ;
        RECT 131.585 23.515 131.755 23.685 ;
        RECT 131.585 18.075 131.755 18.245 ;
        RECT 131.585 12.635 131.755 12.805 ;
        RECT 132.045 56.155 132.215 56.325 ;
        RECT 132.045 50.715 132.215 50.885 ;
        RECT 132.045 45.275 132.215 45.445 ;
        RECT 132.045 39.835 132.215 40.005 ;
        RECT 132.045 34.395 132.215 34.565 ;
        RECT 132.045 28.955 132.215 29.125 ;
        RECT 132.045 23.515 132.215 23.685 ;
        RECT 132.045 18.075 132.215 18.245 ;
        RECT 132.045 12.635 132.215 12.805 ;
        RECT 132.505 56.155 132.675 56.325 ;
        RECT 132.505 50.715 132.675 50.885 ;
        RECT 132.505 45.275 132.675 45.445 ;
        RECT 132.505 39.835 132.675 40.005 ;
        RECT 132.505 34.395 132.675 34.565 ;
        RECT 132.505 28.955 132.675 29.125 ;
        RECT 132.505 23.515 132.675 23.685 ;
        RECT 132.505 18.075 132.675 18.245 ;
        RECT 132.505 12.635 132.675 12.805 ;
        RECT 132.965 56.155 133.135 56.325 ;
        RECT 132.965 50.715 133.135 50.885 ;
        RECT 132.965 45.275 133.135 45.445 ;
        RECT 132.965 39.835 133.135 40.005 ;
        RECT 132.965 34.395 133.135 34.565 ;
        RECT 132.965 28.955 133.135 29.125 ;
        RECT 132.965 23.515 133.135 23.685 ;
        RECT 132.965 18.075 133.135 18.245 ;
        RECT 132.965 12.635 133.135 12.805 ;
        RECT 133.425 56.155 133.595 56.325 ;
        RECT 133.425 50.715 133.595 50.885 ;
        RECT 133.425 45.275 133.595 45.445 ;
        RECT 133.425 39.835 133.595 40.005 ;
        RECT 133.425 34.395 133.595 34.565 ;
        RECT 133.425 28.955 133.595 29.125 ;
        RECT 133.425 23.515 133.595 23.685 ;
        RECT 133.425 18.075 133.595 18.245 ;
        RECT 133.425 12.635 133.595 12.805 ;
        RECT 133.885 56.155 134.055 56.325 ;
        RECT 133.885 50.715 134.055 50.885 ;
        RECT 133.885 45.275 134.055 45.445 ;
        RECT 133.885 39.835 134.055 40.005 ;
        RECT 133.885 34.395 134.055 34.565 ;
        RECT 133.885 28.955 134.055 29.125 ;
        RECT 133.885 23.515 134.055 23.685 ;
        RECT 133.885 18.075 134.055 18.245 ;
        RECT 133.885 12.635 134.055 12.805 ;
        RECT 134.345 56.155 134.515 56.325 ;
        RECT 134.345 50.715 134.515 50.885 ;
        RECT 134.345 45.275 134.515 45.445 ;
        RECT 134.345 39.835 134.515 40.005 ;
        RECT 134.345 34.395 134.515 34.565 ;
        RECT 134.345 28.955 134.515 29.125 ;
        RECT 134.345 23.515 134.515 23.685 ;
        RECT 134.345 18.075 134.515 18.245 ;
        RECT 134.345 12.635 134.515 12.805 ;
        RECT 134.805 56.155 134.975 56.325 ;
        RECT 134.805 50.715 134.975 50.885 ;
        RECT 134.805 45.275 134.975 45.445 ;
        RECT 134.805 39.835 134.975 40.005 ;
        RECT 134.805 34.395 134.975 34.565 ;
        RECT 134.805 28.955 134.975 29.125 ;
        RECT 134.805 23.515 134.975 23.685 ;
        RECT 134.805 18.075 134.975 18.245 ;
        RECT 134.805 12.635 134.975 12.805 ;
        RECT 135.265 56.155 135.435 56.325 ;
        RECT 135.265 50.715 135.435 50.885 ;
        RECT 135.265 45.275 135.435 45.445 ;
        RECT 135.265 39.835 135.435 40.005 ;
        RECT 135.265 34.395 135.435 34.565 ;
        RECT 135.265 28.955 135.435 29.125 ;
        RECT 135.265 23.515 135.435 23.685 ;
        RECT 135.265 18.075 135.435 18.245 ;
        RECT 135.265 12.635 135.435 12.805 ;
        RECT 135.725 56.155 135.895 56.325 ;
        RECT 135.725 50.715 135.895 50.885 ;
        RECT 135.725 45.275 135.895 45.445 ;
        RECT 135.725 39.835 135.895 40.005 ;
        RECT 135.725 34.395 135.895 34.565 ;
        RECT 135.725 28.955 135.895 29.125 ;
        RECT 135.725 23.515 135.895 23.685 ;
        RECT 135.725 18.075 135.895 18.245 ;
        RECT 135.725 12.635 135.895 12.805 ;
        RECT 136.185 56.155 136.355 56.325 ;
        RECT 136.185 50.715 136.355 50.885 ;
        RECT 136.185 45.275 136.355 45.445 ;
        RECT 136.185 39.835 136.355 40.005 ;
        RECT 136.185 34.395 136.355 34.565 ;
        RECT 136.185 28.955 136.355 29.125 ;
        RECT 136.185 23.515 136.355 23.685 ;
        RECT 136.185 18.075 136.355 18.245 ;
        RECT 136.185 12.635 136.355 12.805 ;
        RECT 136.645 56.155 136.815 56.325 ;
        RECT 136.645 50.715 136.815 50.885 ;
        RECT 136.645 45.275 136.815 45.445 ;
        RECT 136.645 39.835 136.815 40.005 ;
        RECT 136.645 34.395 136.815 34.565 ;
        RECT 136.645 28.955 136.815 29.125 ;
        RECT 136.645 23.515 136.815 23.685 ;
        RECT 136.645 18.075 136.815 18.245 ;
        RECT 136.645 12.635 136.815 12.805 ;
        RECT 137.105 56.155 137.275 56.325 ;
        RECT 137.105 50.715 137.275 50.885 ;
        RECT 137.105 45.275 137.275 45.445 ;
        RECT 137.105 39.835 137.275 40.005 ;
        RECT 137.105 34.395 137.275 34.565 ;
        RECT 137.105 28.955 137.275 29.125 ;
        RECT 137.105 23.515 137.275 23.685 ;
        RECT 137.105 18.075 137.275 18.245 ;
        RECT 137.105 12.635 137.275 12.805 ;
        RECT 137.565 56.155 137.735 56.325 ;
        RECT 137.565 50.715 137.735 50.885 ;
        RECT 137.565 45.275 137.735 45.445 ;
        RECT 137.565 39.835 137.735 40.005 ;
        RECT 137.565 34.395 137.735 34.565 ;
        RECT 137.565 28.955 137.735 29.125 ;
        RECT 137.565 23.515 137.735 23.685 ;
        RECT 137.565 18.075 137.735 18.245 ;
        RECT 137.565 12.635 137.735 12.805 ;
        RECT 138.025 56.155 138.195 56.325 ;
        RECT 138.025 50.715 138.195 50.885 ;
        RECT 138.025 45.275 138.195 45.445 ;
        RECT 138.025 39.835 138.195 40.005 ;
        RECT 138.025 34.395 138.195 34.565 ;
        RECT 138.025 28.955 138.195 29.125 ;
        RECT 138.025 23.515 138.195 23.685 ;
        RECT 138.025 18.075 138.195 18.245 ;
        RECT 138.025 12.635 138.195 12.805 ;
        RECT 138.485 56.155 138.655 56.325 ;
        RECT 138.485 50.715 138.655 50.885 ;
        RECT 138.485 45.275 138.655 45.445 ;
        RECT 138.485 39.835 138.655 40.005 ;
        RECT 138.485 34.395 138.655 34.565 ;
        RECT 138.485 28.955 138.655 29.125 ;
        RECT 138.485 23.515 138.655 23.685 ;
        RECT 138.485 18.075 138.655 18.245 ;
        RECT 138.485 12.635 138.655 12.805 ;
        RECT 138.945 56.155 139.115 56.325 ;
        RECT 138.945 50.715 139.115 50.885 ;
        RECT 138.945 45.275 139.115 45.445 ;
        RECT 138.945 39.835 139.115 40.005 ;
        RECT 138.945 34.395 139.115 34.565 ;
        RECT 138.945 28.955 139.115 29.125 ;
        RECT 138.945 23.515 139.115 23.685 ;
        RECT 138.945 18.075 139.115 18.245 ;
        RECT 138.945 12.635 139.115 12.805 ;
        RECT 139.405 56.155 139.575 56.325 ;
        RECT 139.405 50.715 139.575 50.885 ;
        RECT 139.405 45.275 139.575 45.445 ;
        RECT 139.405 39.835 139.575 40.005 ;
        RECT 139.405 34.395 139.575 34.565 ;
        RECT 139.405 28.955 139.575 29.125 ;
        RECT 139.405 23.515 139.575 23.685 ;
        RECT 139.405 18.075 139.575 18.245 ;
        RECT 139.405 12.635 139.575 12.805 ;
        RECT 139.865 56.155 140.035 56.325 ;
        RECT 139.865 50.715 140.035 50.885 ;
        RECT 139.865 45.275 140.035 45.445 ;
        RECT 139.865 39.835 140.035 40.005 ;
        RECT 139.865 34.395 140.035 34.565 ;
        RECT 139.865 28.955 140.035 29.125 ;
        RECT 139.865 23.515 140.035 23.685 ;
        RECT 139.865 18.075 140.035 18.245 ;
        RECT 139.865 12.635 140.035 12.805 ;
        RECT 140.325 56.155 140.495 56.325 ;
        RECT 140.325 50.715 140.495 50.885 ;
        RECT 140.325 45.275 140.495 45.445 ;
        RECT 140.325 39.835 140.495 40.005 ;
        RECT 140.325 34.395 140.495 34.565 ;
        RECT 140.325 28.955 140.495 29.125 ;
        RECT 140.325 23.515 140.495 23.685 ;
        RECT 140.325 18.075 140.495 18.245 ;
        RECT 140.325 12.635 140.495 12.805 ;
        RECT 140.785 56.155 140.955 56.325 ;
        RECT 140.785 50.715 140.955 50.885 ;
        RECT 140.785 45.275 140.955 45.445 ;
        RECT 140.785 39.835 140.955 40.005 ;
        RECT 140.785 34.395 140.955 34.565 ;
        RECT 140.785 28.955 140.955 29.125 ;
        RECT 140.785 23.515 140.955 23.685 ;
        RECT 140.785 18.075 140.955 18.245 ;
        RECT 140.785 12.635 140.955 12.805 ;
        RECT 141.245 56.155 141.415 56.325 ;
        RECT 141.245 50.715 141.415 50.885 ;
        RECT 141.245 45.275 141.415 45.445 ;
        RECT 141.245 39.835 141.415 40.005 ;
        RECT 141.245 34.395 141.415 34.565 ;
        RECT 141.245 28.955 141.415 29.125 ;
        RECT 141.245 23.515 141.415 23.685 ;
        RECT 141.245 18.075 141.415 18.245 ;
        RECT 141.245 12.635 141.415 12.805 ;
        RECT 141.705 56.155 141.875 56.325 ;
        RECT 141.705 50.715 141.875 50.885 ;
        RECT 141.705 45.275 141.875 45.445 ;
        RECT 141.705 39.835 141.875 40.005 ;
        RECT 141.705 34.395 141.875 34.565 ;
        RECT 141.705 28.955 141.875 29.125 ;
        RECT 141.705 23.515 141.875 23.685 ;
        RECT 141.705 18.075 141.875 18.245 ;
        RECT 141.705 12.635 141.875 12.805 ;
        RECT 142.165 56.155 142.335 56.325 ;
        RECT 142.165 50.715 142.335 50.885 ;
        RECT 142.165 45.275 142.335 45.445 ;
        RECT 142.165 39.835 142.335 40.005 ;
        RECT 142.165 34.395 142.335 34.565 ;
        RECT 142.165 28.955 142.335 29.125 ;
        RECT 142.165 23.515 142.335 23.685 ;
        RECT 142.165 18.075 142.335 18.245 ;
        RECT 142.165 12.635 142.335 12.805 ;
        RECT 142.625 56.155 142.795 56.325 ;
        RECT 142.625 50.715 142.795 50.885 ;
        RECT 142.625 45.275 142.795 45.445 ;
        RECT 142.625 39.835 142.795 40.005 ;
        RECT 142.625 34.395 142.795 34.565 ;
        RECT 142.625 28.955 142.795 29.125 ;
        RECT 142.625 23.515 142.795 23.685 ;
        RECT 142.625 18.075 142.795 18.245 ;
        RECT 142.625 12.635 142.795 12.805 ;
        RECT 143.085 56.155 143.255 56.325 ;
        RECT 143.085 50.715 143.255 50.885 ;
        RECT 143.085 45.275 143.255 45.445 ;
        RECT 143.085 39.835 143.255 40.005 ;
        RECT 143.085 34.395 143.255 34.565 ;
        RECT 143.085 28.955 143.255 29.125 ;
        RECT 143.085 23.515 143.255 23.685 ;
        RECT 143.085 18.075 143.255 18.245 ;
        RECT 143.085 12.635 143.255 12.805 ;
        RECT 143.545 56.155 143.715 56.325 ;
        RECT 143.545 50.715 143.715 50.885 ;
        RECT 143.545 45.275 143.715 45.445 ;
        RECT 143.545 39.835 143.715 40.005 ;
        RECT 143.545 34.395 143.715 34.565 ;
        RECT 143.545 28.955 143.715 29.125 ;
        RECT 143.545 23.515 143.715 23.685 ;
        RECT 143.545 18.075 143.715 18.245 ;
        RECT 143.545 12.635 143.715 12.805 ;
        RECT 144.005 56.155 144.175 56.325 ;
        RECT 144.005 50.715 144.175 50.885 ;
        RECT 144.005 45.275 144.175 45.445 ;
        RECT 144.005 39.835 144.175 40.005 ;
        RECT 144.005 34.395 144.175 34.565 ;
        RECT 144.005 28.955 144.175 29.125 ;
        RECT 144.005 23.515 144.175 23.685 ;
        RECT 144.005 18.075 144.175 18.245 ;
        RECT 144.005 12.635 144.175 12.805 ;
        RECT 144.465 56.155 144.635 56.325 ;
        RECT 144.465 50.715 144.635 50.885 ;
        RECT 144.465 45.275 144.635 45.445 ;
        RECT 144.465 39.835 144.635 40.005 ;
        RECT 144.465 34.395 144.635 34.565 ;
        RECT 144.465 28.955 144.635 29.125 ;
        RECT 144.465 23.515 144.635 23.685 ;
        RECT 144.465 18.075 144.635 18.245 ;
        RECT 144.465 12.635 144.635 12.805 ;
        RECT 144.925 56.155 145.095 56.325 ;
        RECT 144.925 50.715 145.095 50.885 ;
        RECT 144.925 45.275 145.095 45.445 ;
        RECT 144.925 39.835 145.095 40.005 ;
        RECT 144.925 34.395 145.095 34.565 ;
        RECT 144.925 28.955 145.095 29.125 ;
        RECT 144.925 23.515 145.095 23.685 ;
        RECT 144.925 18.075 145.095 18.245 ;
        RECT 144.925 12.635 145.095 12.805 ;
        RECT 145.385 56.155 145.555 56.325 ;
        RECT 145.385 50.715 145.555 50.885 ;
        RECT 145.385 45.275 145.555 45.445 ;
        RECT 145.385 39.835 145.555 40.005 ;
        RECT 145.385 34.395 145.555 34.565 ;
        RECT 145.385 28.955 145.555 29.125 ;
        RECT 145.385 23.515 145.555 23.685 ;
        RECT 145.385 18.075 145.555 18.245 ;
        RECT 145.385 12.635 145.555 12.805 ;
        RECT 145.845 56.155 146.015 56.325 ;
        RECT 145.845 50.715 146.015 50.885 ;
        RECT 145.845 45.275 146.015 45.445 ;
        RECT 145.845 39.835 146.015 40.005 ;
        RECT 145.845 34.395 146.015 34.565 ;
        RECT 145.845 28.955 146.015 29.125 ;
        RECT 145.845 23.515 146.015 23.685 ;
        RECT 145.845 18.075 146.015 18.245 ;
        RECT 145.845 12.635 146.015 12.805 ;
        RECT 146.305 56.155 146.475 56.325 ;
        RECT 146.305 50.715 146.475 50.885 ;
        RECT 146.305 45.275 146.475 45.445 ;
        RECT 146.305 39.835 146.475 40.005 ;
        RECT 146.305 34.395 146.475 34.565 ;
        RECT 146.305 28.955 146.475 29.125 ;
        RECT 146.305 23.515 146.475 23.685 ;
        RECT 146.305 18.075 146.475 18.245 ;
        RECT 146.305 12.635 146.475 12.805 ;
        RECT 146.765 56.155 146.935 56.325 ;
        RECT 146.765 50.715 146.935 50.885 ;
        RECT 146.765 45.275 146.935 45.445 ;
        RECT 146.765 39.835 146.935 40.005 ;
        RECT 146.765 34.395 146.935 34.565 ;
        RECT 146.765 28.955 146.935 29.125 ;
        RECT 146.765 23.515 146.935 23.685 ;
        RECT 146.765 18.075 146.935 18.245 ;
        RECT 146.765 12.635 146.935 12.805 ;
        RECT 147.225 56.155 147.395 56.325 ;
        RECT 147.225 50.715 147.395 50.885 ;
        RECT 147.225 45.275 147.395 45.445 ;
        RECT 147.225 39.835 147.395 40.005 ;
        RECT 147.225 34.395 147.395 34.565 ;
        RECT 147.225 28.955 147.395 29.125 ;
        RECT 147.225 23.515 147.395 23.685 ;
        RECT 147.225 18.075 147.395 18.245 ;
        RECT 147.225 12.635 147.395 12.805 ;
        RECT 147.685 56.155 147.855 56.325 ;
        RECT 147.685 50.715 147.855 50.885 ;
        RECT 147.685 45.275 147.855 45.445 ;
        RECT 147.685 39.835 147.855 40.005 ;
        RECT 147.685 34.395 147.855 34.565 ;
        RECT 147.685 28.955 147.855 29.125 ;
        RECT 147.685 23.515 147.855 23.685 ;
        RECT 147.685 18.075 147.855 18.245 ;
        RECT 147.685 12.635 147.855 12.805 ;
        RECT 148.145 56.155 148.315 56.325 ;
        RECT 148.145 50.715 148.315 50.885 ;
        RECT 148.145 45.275 148.315 45.445 ;
        RECT 148.145 39.835 148.315 40.005 ;
        RECT 148.145 34.395 148.315 34.565 ;
        RECT 148.145 28.955 148.315 29.125 ;
        RECT 148.145 23.515 148.315 23.685 ;
        RECT 148.145 18.075 148.315 18.245 ;
        RECT 148.145 12.635 148.315 12.805 ;
        RECT 148.605 56.155 148.775 56.325 ;
        RECT 148.605 50.715 148.775 50.885 ;
        RECT 148.605 45.275 148.775 45.445 ;
        RECT 148.605 39.835 148.775 40.005 ;
        RECT 148.605 34.395 148.775 34.565 ;
        RECT 148.605 28.955 148.775 29.125 ;
        RECT 148.605 23.515 148.775 23.685 ;
        RECT 148.605 18.075 148.775 18.245 ;
        RECT 148.605 12.635 148.775 12.805 ;
        RECT 149.065 56.155 149.235 56.325 ;
        RECT 149.065 50.715 149.235 50.885 ;
        RECT 149.065 45.275 149.235 45.445 ;
        RECT 149.065 39.835 149.235 40.005 ;
        RECT 149.065 34.395 149.235 34.565 ;
        RECT 149.065 28.955 149.235 29.125 ;
        RECT 149.065 23.515 149.235 23.685 ;
        RECT 149.065 18.075 149.235 18.245 ;
        RECT 149.065 12.635 149.235 12.805 ;
        RECT 149.525 56.155 149.695 56.325 ;
        RECT 149.525 50.715 149.695 50.885 ;
        RECT 149.525 45.275 149.695 45.445 ;
        RECT 149.525 39.835 149.695 40.005 ;
        RECT 149.525 34.395 149.695 34.565 ;
        RECT 149.525 28.955 149.695 29.125 ;
        RECT 149.525 23.515 149.695 23.685 ;
        RECT 149.525 18.075 149.695 18.245 ;
        RECT 149.525 12.635 149.695 12.805 ;
        RECT 149.985 56.155 150.155 56.325 ;
        RECT 149.985 50.715 150.155 50.885 ;
        RECT 149.985 45.275 150.155 45.445 ;
        RECT 149.985 39.835 150.155 40.005 ;
        RECT 149.985 34.395 150.155 34.565 ;
        RECT 149.985 28.955 150.155 29.125 ;
        RECT 149.985 23.515 150.155 23.685 ;
        RECT 149.985 18.075 150.155 18.245 ;
        RECT 149.985 12.635 150.155 12.805 ;
        RECT 150.445 56.155 150.615 56.325 ;
        RECT 150.445 50.715 150.615 50.885 ;
        RECT 150.445 45.275 150.615 45.445 ;
        RECT 150.445 39.835 150.615 40.005 ;
        RECT 150.445 34.395 150.615 34.565 ;
        RECT 150.445 28.955 150.615 29.125 ;
        RECT 150.445 23.515 150.615 23.685 ;
        RECT 150.445 18.075 150.615 18.245 ;
        RECT 150.445 12.635 150.615 12.805 ;
        RECT 150.905 56.155 151.075 56.325 ;
        RECT 150.905 50.715 151.075 50.885 ;
        RECT 150.905 45.275 151.075 45.445 ;
        RECT 150.905 39.835 151.075 40.005 ;
        RECT 150.905 34.395 151.075 34.565 ;
        RECT 150.905 28.955 151.075 29.125 ;
        RECT 150.905 23.515 151.075 23.685 ;
        RECT 150.905 18.075 151.075 18.245 ;
        RECT 150.905 12.635 151.075 12.805 ;
        RECT 151.365 56.155 151.535 56.325 ;
        RECT 151.365 50.715 151.535 50.885 ;
        RECT 151.365 45.275 151.535 45.445 ;
        RECT 151.365 39.835 151.535 40.005 ;
        RECT 151.365 34.395 151.535 34.565 ;
        RECT 151.365 28.955 151.535 29.125 ;
        RECT 151.365 23.515 151.535 23.685 ;
        RECT 151.365 18.075 151.535 18.245 ;
        RECT 151.365 12.635 151.535 12.805 ;
        RECT 151.825 56.155 151.995 56.325 ;
        RECT 151.825 50.715 151.995 50.885 ;
        RECT 151.825 45.275 151.995 45.445 ;
        RECT 151.825 39.835 151.995 40.005 ;
        RECT 151.825 34.395 151.995 34.565 ;
        RECT 151.825 28.955 151.995 29.125 ;
        RECT 151.825 23.515 151.995 23.685 ;
        RECT 151.825 18.075 151.995 18.245 ;
        RECT 151.825 12.635 151.995 12.805 ;
        RECT 152.285 56.155 152.455 56.325 ;
        RECT 152.285 50.715 152.455 50.885 ;
        RECT 152.285 45.275 152.455 45.445 ;
        RECT 152.285 39.835 152.455 40.005 ;
        RECT 152.285 34.395 152.455 34.565 ;
        RECT 152.285 28.955 152.455 29.125 ;
        RECT 152.285 23.515 152.455 23.685 ;
        RECT 152.285 18.075 152.455 18.245 ;
        RECT 152.285 12.635 152.455 12.805 ;
        RECT 152.745 56.155 152.915 56.325 ;
        RECT 152.745 50.715 152.915 50.885 ;
        RECT 152.745 45.275 152.915 45.445 ;
        RECT 152.745 39.835 152.915 40.005 ;
        RECT 152.745 34.395 152.915 34.565 ;
        RECT 152.745 28.955 152.915 29.125 ;
        RECT 152.745 23.515 152.915 23.685 ;
        RECT 152.745 18.075 152.915 18.245 ;
        RECT 152.745 12.635 152.915 12.805 ;
        RECT 153.205 56.155 153.375 56.325 ;
        RECT 153.205 50.715 153.375 50.885 ;
        RECT 153.205 45.275 153.375 45.445 ;
        RECT 153.205 39.835 153.375 40.005 ;
        RECT 153.205 34.395 153.375 34.565 ;
        RECT 153.205 28.955 153.375 29.125 ;
        RECT 153.205 23.515 153.375 23.685 ;
        RECT 153.205 18.075 153.375 18.245 ;
        RECT 153.205 12.635 153.375 12.805 ;
        RECT 153.665 56.155 153.835 56.325 ;
        RECT 153.665 50.715 153.835 50.885 ;
        RECT 153.665 45.275 153.835 45.445 ;
        RECT 153.665 39.835 153.835 40.005 ;
        RECT 153.665 34.395 153.835 34.565 ;
        RECT 153.665 28.955 153.835 29.125 ;
        RECT 153.665 23.515 153.835 23.685 ;
        RECT 153.665 18.075 153.835 18.245 ;
        RECT 153.665 12.635 153.835 12.805 ;
        RECT 154.125 56.155 154.295 56.325 ;
        RECT 154.125 50.715 154.295 50.885 ;
        RECT 154.125 45.275 154.295 45.445 ;
        RECT 154.125 39.835 154.295 40.005 ;
        RECT 154.125 34.395 154.295 34.565 ;
        RECT 154.125 28.955 154.295 29.125 ;
        RECT 154.125 23.515 154.295 23.685 ;
        RECT 154.125 18.075 154.295 18.245 ;
        RECT 154.125 12.635 154.295 12.805 ;
        RECT 154.585 56.155 154.755 56.325 ;
        RECT 154.585 50.715 154.755 50.885 ;
        RECT 154.585 45.275 154.755 45.445 ;
        RECT 154.585 39.835 154.755 40.005 ;
        RECT 154.585 34.395 154.755 34.565 ;
        RECT 154.585 28.955 154.755 29.125 ;
        RECT 154.585 23.515 154.755 23.685 ;
        RECT 154.585 18.075 154.755 18.245 ;
        RECT 154.585 12.635 154.755 12.805 ;
        RECT 155.045 56.155 155.215 56.325 ;
        RECT 155.045 50.715 155.215 50.885 ;
        RECT 155.045 45.275 155.215 45.445 ;
        RECT 155.045 39.835 155.215 40.005 ;
        RECT 155.045 34.395 155.215 34.565 ;
        RECT 155.045 28.955 155.215 29.125 ;
        RECT 155.045 23.515 155.215 23.685 ;
        RECT 155.045 18.075 155.215 18.245 ;
        RECT 155.045 12.635 155.215 12.805 ;
        RECT 155.505 56.155 155.675 56.325 ;
        RECT 155.505 50.715 155.675 50.885 ;
        RECT 155.505 45.275 155.675 45.445 ;
        RECT 155.505 39.835 155.675 40.005 ;
        RECT 155.505 34.395 155.675 34.565 ;
        RECT 155.505 28.955 155.675 29.125 ;
        RECT 155.505 23.515 155.675 23.685 ;
        RECT 155.505 18.075 155.675 18.245 ;
        RECT 155.505 12.635 155.675 12.805 ;
        RECT 155.965 56.155 156.135 56.325 ;
        RECT 155.965 50.715 156.135 50.885 ;
        RECT 155.965 45.275 156.135 45.445 ;
        RECT 155.965 39.835 156.135 40.005 ;
        RECT 155.965 34.395 156.135 34.565 ;
        RECT 155.965 28.955 156.135 29.125 ;
        RECT 155.965 23.515 156.135 23.685 ;
        RECT 155.965 18.075 156.135 18.245 ;
        RECT 155.965 12.635 156.135 12.805 ;
        RECT 156.425 56.155 156.595 56.325 ;
        RECT 156.425 50.715 156.595 50.885 ;
        RECT 156.425 45.275 156.595 45.445 ;
        RECT 156.425 39.835 156.595 40.005 ;
        RECT 156.425 34.395 156.595 34.565 ;
        RECT 156.425 28.955 156.595 29.125 ;
        RECT 156.425 23.515 156.595 23.685 ;
        RECT 156.425 18.075 156.595 18.245 ;
        RECT 156.425 12.635 156.595 12.805 ;
        RECT 156.885 56.155 157.055 56.325 ;
        RECT 156.885 50.715 157.055 50.885 ;
        RECT 156.885 45.275 157.055 45.445 ;
        RECT 156.885 39.835 157.055 40.005 ;
        RECT 156.885 34.395 157.055 34.565 ;
        RECT 156.885 28.955 157.055 29.125 ;
        RECT 156.885 23.515 157.055 23.685 ;
        RECT 156.885 18.075 157.055 18.245 ;
        RECT 156.885 12.635 157.055 12.805 ;
        RECT 157.345 56.155 157.515 56.325 ;
        RECT 157.345 50.715 157.515 50.885 ;
        RECT 157.345 45.275 157.515 45.445 ;
        RECT 157.345 39.835 157.515 40.005 ;
        RECT 157.345 34.395 157.515 34.565 ;
        RECT 157.345 28.955 157.515 29.125 ;
        RECT 157.345 23.515 157.515 23.685 ;
        RECT 157.345 18.075 157.515 18.245 ;
        RECT 157.345 12.635 157.515 12.805 ;
        RECT 157.805 56.155 157.975 56.325 ;
        RECT 157.805 50.715 157.975 50.885 ;
        RECT 157.805 45.275 157.975 45.445 ;
        RECT 157.805 39.835 157.975 40.005 ;
        RECT 157.805 34.395 157.975 34.565 ;
        RECT 157.805 28.955 157.975 29.125 ;
        RECT 157.805 23.515 157.975 23.685 ;
        RECT 157.805 18.075 157.975 18.245 ;
        RECT 157.805 12.635 157.975 12.805 ;
        RECT 158.265 56.155 158.435 56.325 ;
        RECT 158.265 50.715 158.435 50.885 ;
        RECT 158.265 45.275 158.435 45.445 ;
        RECT 158.265 39.835 158.435 40.005 ;
        RECT 158.265 34.395 158.435 34.565 ;
        RECT 158.265 28.955 158.435 29.125 ;
        RECT 158.265 23.515 158.435 23.685 ;
        RECT 158.265 18.075 158.435 18.245 ;
        RECT 158.265 12.635 158.435 12.805 ;
        RECT 158.725 56.155 158.895 56.325 ;
        RECT 158.725 50.715 158.895 50.885 ;
        RECT 158.725 45.275 158.895 45.445 ;
        RECT 158.725 39.835 158.895 40.005 ;
        RECT 158.725 34.395 158.895 34.565 ;
        RECT 158.725 28.955 158.895 29.125 ;
        RECT 158.725 23.515 158.895 23.685 ;
        RECT 158.725 18.075 158.895 18.245 ;
        RECT 158.725 12.635 158.895 12.805 ;
        RECT 159.185 56.155 159.355 56.325 ;
        RECT 159.185 50.715 159.355 50.885 ;
        RECT 159.185 45.275 159.355 45.445 ;
        RECT 159.185 39.835 159.355 40.005 ;
        RECT 159.185 34.395 159.355 34.565 ;
        RECT 159.185 28.955 159.355 29.125 ;
        RECT 159.185 23.515 159.355 23.685 ;
        RECT 159.185 18.075 159.355 18.245 ;
        RECT 159.185 12.635 159.355 12.805 ;
        RECT 159.645 56.155 159.815 56.325 ;
        RECT 159.645 50.715 159.815 50.885 ;
        RECT 159.645 45.275 159.815 45.445 ;
        RECT 159.645 39.835 159.815 40.005 ;
        RECT 159.645 34.395 159.815 34.565 ;
        RECT 159.645 28.955 159.815 29.125 ;
        RECT 159.645 23.515 159.815 23.685 ;
        RECT 159.645 18.075 159.815 18.245 ;
        RECT 159.645 12.635 159.815 12.805 ;
        RECT 160.105 56.155 160.275 56.325 ;
        RECT 160.105 50.715 160.275 50.885 ;
        RECT 160.105 45.275 160.275 45.445 ;
        RECT 160.105 39.835 160.275 40.005 ;
        RECT 160.105 34.395 160.275 34.565 ;
        RECT 160.105 28.955 160.275 29.125 ;
        RECT 160.105 23.515 160.275 23.685 ;
        RECT 160.105 18.075 160.275 18.245 ;
        RECT 160.105 12.635 160.275 12.805 ;
        RECT 160.565 56.155 160.735 56.325 ;
        RECT 160.565 50.715 160.735 50.885 ;
        RECT 160.565 45.275 160.735 45.445 ;
        RECT 160.565 39.835 160.735 40.005 ;
        RECT 160.565 34.395 160.735 34.565 ;
        RECT 160.565 28.955 160.735 29.125 ;
        RECT 160.565 23.515 160.735 23.685 ;
        RECT 160.565 18.075 160.735 18.245 ;
        RECT 160.565 12.635 160.735 12.805 ;
        RECT 161.025 56.155 161.195 56.325 ;
        RECT 161.025 50.715 161.195 50.885 ;
        RECT 161.025 45.275 161.195 45.445 ;
        RECT 161.025 39.835 161.195 40.005 ;
        RECT 161.025 34.395 161.195 34.565 ;
        RECT 161.025 28.955 161.195 29.125 ;
        RECT 161.025 23.515 161.195 23.685 ;
        RECT 161.025 18.075 161.195 18.245 ;
        RECT 161.025 12.635 161.195 12.805 ;
        RECT 161.485 56.155 161.655 56.325 ;
        RECT 161.485 50.715 161.655 50.885 ;
        RECT 161.485 45.275 161.655 45.445 ;
        RECT 161.485 39.835 161.655 40.005 ;
        RECT 161.485 34.395 161.655 34.565 ;
        RECT 161.485 28.955 161.655 29.125 ;
        RECT 161.485 23.515 161.655 23.685 ;
        RECT 161.485 18.075 161.655 18.245 ;
        RECT 161.485 12.635 161.655 12.805 ;
        RECT 161.945 56.155 162.115 56.325 ;
        RECT 161.945 50.715 162.115 50.885 ;
        RECT 161.945 45.275 162.115 45.445 ;
        RECT 161.945 39.835 162.115 40.005 ;
        RECT 161.945 34.395 162.115 34.565 ;
        RECT 161.945 28.955 162.115 29.125 ;
        RECT 161.945 23.515 162.115 23.685 ;
        RECT 161.945 18.075 162.115 18.245 ;
        RECT 161.945 12.635 162.115 12.805 ;
        RECT 162.405 56.155 162.575 56.325 ;
        RECT 162.405 50.715 162.575 50.885 ;
        RECT 162.405 45.275 162.575 45.445 ;
        RECT 162.405 39.835 162.575 40.005 ;
        RECT 162.405 34.395 162.575 34.565 ;
        RECT 162.405 28.955 162.575 29.125 ;
        RECT 162.405 23.515 162.575 23.685 ;
        RECT 162.405 18.075 162.575 18.245 ;
        RECT 162.405 12.635 162.575 12.805 ;
        RECT 162.865 56.155 163.035 56.325 ;
        RECT 162.865 50.715 163.035 50.885 ;
        RECT 162.865 45.275 163.035 45.445 ;
        RECT 162.865 39.835 163.035 40.005 ;
        RECT 162.865 34.395 163.035 34.565 ;
        RECT 162.865 28.955 163.035 29.125 ;
        RECT 162.865 23.515 163.035 23.685 ;
        RECT 162.865 18.075 163.035 18.245 ;
        RECT 162.865 12.635 163.035 12.805 ;
        RECT 163.325 56.155 163.495 56.325 ;
        RECT 163.325 50.715 163.495 50.885 ;
        RECT 163.325 45.275 163.495 45.445 ;
        RECT 61.205 50.715 61.375 50.885 ;
        RECT 61.205 45.275 61.375 45.445 ;
        RECT 61.205 39.835 61.375 40.005 ;
        RECT 61.205 34.395 61.375 34.565 ;
        RECT 61.205 28.955 61.375 29.125 ;
        RECT 61.205 23.515 61.375 23.685 ;
        RECT 61.205 18.075 61.375 18.245 ;
        RECT 61.205 12.635 61.375 12.805 ;
        RECT 61.665 56.155 61.835 56.325 ;
        RECT 61.665 50.715 61.835 50.885 ;
        RECT 61.665 45.275 61.835 45.445 ;
        RECT 61.665 39.835 61.835 40.005 ;
        RECT 61.665 34.395 61.835 34.565 ;
        RECT 61.665 28.955 61.835 29.125 ;
        RECT 61.665 23.515 61.835 23.685 ;
        RECT 61.665 18.075 61.835 18.245 ;
        RECT 61.665 12.635 61.835 12.805 ;
        RECT 62.125 56.155 62.295 56.325 ;
        RECT 62.125 50.715 62.295 50.885 ;
        RECT 62.125 45.275 62.295 45.445 ;
        RECT 62.125 39.835 62.295 40.005 ;
        RECT 62.125 34.395 62.295 34.565 ;
        RECT 62.125 28.955 62.295 29.125 ;
        RECT 62.125 23.515 62.295 23.685 ;
        RECT 62.125 18.075 62.295 18.245 ;
        RECT 62.125 12.635 62.295 12.805 ;
        RECT 62.585 56.155 62.755 56.325 ;
        RECT 62.585 50.715 62.755 50.885 ;
        RECT 62.585 45.275 62.755 45.445 ;
        RECT 62.585 39.835 62.755 40.005 ;
        RECT 62.585 34.395 62.755 34.565 ;
        RECT 62.585 28.955 62.755 29.125 ;
        RECT 62.585 23.515 62.755 23.685 ;
        RECT 62.585 18.075 62.755 18.245 ;
        RECT 62.585 12.635 62.755 12.805 ;
        RECT 63.045 56.155 63.215 56.325 ;
        RECT 63.045 50.715 63.215 50.885 ;
        RECT 63.045 45.275 63.215 45.445 ;
        RECT 63.045 39.835 63.215 40.005 ;
        RECT 63.045 34.395 63.215 34.565 ;
        RECT 63.045 28.955 63.215 29.125 ;
        RECT 63.045 23.515 63.215 23.685 ;
        RECT 63.045 18.075 63.215 18.245 ;
        RECT 63.045 12.635 63.215 12.805 ;
        RECT 63.505 56.155 63.675 56.325 ;
        RECT 63.505 50.715 63.675 50.885 ;
        RECT 63.505 45.275 63.675 45.445 ;
        RECT 63.505 39.835 63.675 40.005 ;
        RECT 63.505 34.395 63.675 34.565 ;
        RECT 63.505 28.955 63.675 29.125 ;
        RECT 63.505 23.515 63.675 23.685 ;
        RECT 63.505 18.075 63.675 18.245 ;
        RECT 63.505 12.635 63.675 12.805 ;
        RECT 63.965 56.155 64.135 56.325 ;
        RECT 63.965 50.715 64.135 50.885 ;
        RECT 63.965 45.275 64.135 45.445 ;
        RECT 63.965 39.835 64.135 40.005 ;
        RECT 63.965 34.395 64.135 34.565 ;
        RECT 63.965 28.955 64.135 29.125 ;
        RECT 63.965 23.515 64.135 23.685 ;
        RECT 63.965 18.075 64.135 18.245 ;
        RECT 63.965 12.635 64.135 12.805 ;
        RECT 64.425 56.155 64.595 56.325 ;
        RECT 64.425 50.715 64.595 50.885 ;
        RECT 64.425 45.275 64.595 45.445 ;
        RECT 64.425 39.835 64.595 40.005 ;
        RECT 64.425 34.395 64.595 34.565 ;
        RECT 64.425 28.955 64.595 29.125 ;
        RECT 64.425 23.515 64.595 23.685 ;
        RECT 64.425 18.075 64.595 18.245 ;
        RECT 64.425 12.635 64.595 12.805 ;
        RECT 64.885 56.155 65.055 56.325 ;
        RECT 64.885 50.715 65.055 50.885 ;
        RECT 64.885 45.275 65.055 45.445 ;
        RECT 64.885 39.835 65.055 40.005 ;
        RECT 64.885 34.395 65.055 34.565 ;
        RECT 64.885 28.955 65.055 29.125 ;
        RECT 64.885 23.515 65.055 23.685 ;
        RECT 64.885 18.075 65.055 18.245 ;
        RECT 64.885 12.635 65.055 12.805 ;
        RECT 65.345 56.155 65.515 56.325 ;
        RECT 65.345 50.715 65.515 50.885 ;
        RECT 65.345 45.275 65.515 45.445 ;
        RECT 65.345 39.835 65.515 40.005 ;
        RECT 65.345 34.395 65.515 34.565 ;
        RECT 65.345 28.955 65.515 29.125 ;
        RECT 65.345 23.515 65.515 23.685 ;
        RECT 65.345 18.075 65.515 18.245 ;
        RECT 65.345 12.635 65.515 12.805 ;
        RECT 65.805 56.155 65.975 56.325 ;
        RECT 65.805 50.715 65.975 50.885 ;
        RECT 65.805 45.275 65.975 45.445 ;
        RECT 65.805 39.835 65.975 40.005 ;
        RECT 65.805 34.395 65.975 34.565 ;
        RECT 65.805 28.955 65.975 29.125 ;
        RECT 65.805 23.515 65.975 23.685 ;
        RECT 65.805 18.075 65.975 18.245 ;
        RECT 65.805 12.635 65.975 12.805 ;
        RECT 66.265 56.155 66.435 56.325 ;
        RECT 66.265 50.715 66.435 50.885 ;
        RECT 66.265 45.275 66.435 45.445 ;
        RECT 66.265 39.835 66.435 40.005 ;
        RECT 66.265 34.395 66.435 34.565 ;
        RECT 66.265 28.955 66.435 29.125 ;
        RECT 66.265 23.515 66.435 23.685 ;
        RECT 66.265 18.075 66.435 18.245 ;
        RECT 66.265 12.635 66.435 12.805 ;
        RECT 66.725 56.155 66.895 56.325 ;
        RECT 66.725 50.715 66.895 50.885 ;
        RECT 66.725 45.275 66.895 45.445 ;
        RECT 66.725 39.835 66.895 40.005 ;
        RECT 66.725 34.395 66.895 34.565 ;
        RECT 66.725 28.955 66.895 29.125 ;
        RECT 66.725 23.515 66.895 23.685 ;
        RECT 66.725 18.075 66.895 18.245 ;
        RECT 66.725 12.635 66.895 12.805 ;
        RECT 67.185 56.155 67.355 56.325 ;
        RECT 67.185 50.715 67.355 50.885 ;
        RECT 67.185 45.275 67.355 45.445 ;
        RECT 67.185 39.835 67.355 40.005 ;
        RECT 67.185 34.395 67.355 34.565 ;
        RECT 67.185 28.955 67.355 29.125 ;
        RECT 67.185 23.515 67.355 23.685 ;
        RECT 67.185 18.075 67.355 18.245 ;
        RECT 67.185 12.635 67.355 12.805 ;
        RECT 67.645 56.155 67.815 56.325 ;
        RECT 67.645 50.715 67.815 50.885 ;
        RECT 67.645 45.275 67.815 45.445 ;
        RECT 67.645 39.835 67.815 40.005 ;
        RECT 67.645 34.395 67.815 34.565 ;
        RECT 67.645 28.955 67.815 29.125 ;
        RECT 67.645 23.515 67.815 23.685 ;
        RECT 67.645 18.075 67.815 18.245 ;
        RECT 67.645 12.635 67.815 12.805 ;
        RECT 68.105 56.155 68.275 56.325 ;
        RECT 68.105 50.715 68.275 50.885 ;
        RECT 68.105 45.275 68.275 45.445 ;
        RECT 68.105 39.835 68.275 40.005 ;
        RECT 68.105 34.395 68.275 34.565 ;
        RECT 68.105 28.955 68.275 29.125 ;
        RECT 68.105 23.515 68.275 23.685 ;
        RECT 68.105 18.075 68.275 18.245 ;
        RECT 68.105 12.635 68.275 12.805 ;
        RECT 68.565 56.155 68.735 56.325 ;
        RECT 68.565 50.715 68.735 50.885 ;
        RECT 68.565 45.275 68.735 45.445 ;
        RECT 68.565 39.835 68.735 40.005 ;
        RECT 68.565 34.395 68.735 34.565 ;
        RECT 68.565 28.955 68.735 29.125 ;
        RECT 68.565 23.515 68.735 23.685 ;
        RECT 68.565 18.075 68.735 18.245 ;
        RECT 68.565 12.635 68.735 12.805 ;
        RECT 69.025 56.155 69.195 56.325 ;
        RECT 69.025 50.715 69.195 50.885 ;
        RECT 69.025 45.275 69.195 45.445 ;
        RECT 69.025 39.835 69.195 40.005 ;
        RECT 69.025 34.395 69.195 34.565 ;
        RECT 69.025 28.955 69.195 29.125 ;
        RECT 69.025 23.515 69.195 23.685 ;
        RECT 69.025 18.075 69.195 18.245 ;
        RECT 69.025 12.635 69.195 12.805 ;
        RECT 69.485 56.155 69.655 56.325 ;
        RECT 69.485 50.715 69.655 50.885 ;
        RECT 69.485 45.275 69.655 45.445 ;
        RECT 69.485 39.835 69.655 40.005 ;
        RECT 69.485 34.395 69.655 34.565 ;
        RECT 69.485 28.955 69.655 29.125 ;
        RECT 69.485 23.515 69.655 23.685 ;
        RECT 69.485 18.075 69.655 18.245 ;
        RECT 69.485 12.635 69.655 12.805 ;
        RECT 69.945 56.155 70.115 56.325 ;
        RECT 69.945 50.715 70.115 50.885 ;
        RECT 69.945 45.275 70.115 45.445 ;
        RECT 69.945 39.835 70.115 40.005 ;
        RECT 69.945 34.395 70.115 34.565 ;
        RECT 69.945 28.955 70.115 29.125 ;
        RECT 69.945 23.515 70.115 23.685 ;
        RECT 69.945 18.075 70.115 18.245 ;
        RECT 69.945 12.635 70.115 12.805 ;
        RECT 70.405 56.155 70.575 56.325 ;
        RECT 70.405 50.715 70.575 50.885 ;
        RECT 70.405 45.275 70.575 45.445 ;
        RECT 70.405 39.835 70.575 40.005 ;
        RECT 70.405 34.395 70.575 34.565 ;
        RECT 70.405 28.955 70.575 29.125 ;
        RECT 70.405 23.515 70.575 23.685 ;
        RECT 70.405 18.075 70.575 18.245 ;
        RECT 70.405 12.635 70.575 12.805 ;
        RECT 70.865 56.155 71.035 56.325 ;
        RECT 70.865 50.715 71.035 50.885 ;
        RECT 70.865 45.275 71.035 45.445 ;
        RECT 70.865 39.835 71.035 40.005 ;
        RECT 70.865 34.395 71.035 34.565 ;
        RECT 70.865 28.955 71.035 29.125 ;
        RECT 70.865 23.515 71.035 23.685 ;
        RECT 70.865 18.075 71.035 18.245 ;
        RECT 70.865 12.635 71.035 12.805 ;
        RECT 71.325 56.155 71.495 56.325 ;
        RECT 71.325 50.715 71.495 50.885 ;
        RECT 71.325 45.275 71.495 45.445 ;
        RECT 71.325 39.835 71.495 40.005 ;
        RECT 71.325 34.395 71.495 34.565 ;
        RECT 71.325 28.955 71.495 29.125 ;
        RECT 71.325 23.515 71.495 23.685 ;
        RECT 71.325 18.075 71.495 18.245 ;
        RECT 71.325 12.635 71.495 12.805 ;
        RECT 71.785 56.155 71.955 56.325 ;
        RECT 71.785 50.715 71.955 50.885 ;
        RECT 71.785 45.275 71.955 45.445 ;
        RECT 71.785 39.835 71.955 40.005 ;
        RECT 71.785 34.395 71.955 34.565 ;
        RECT 71.785 28.955 71.955 29.125 ;
        RECT 71.785 23.515 71.955 23.685 ;
        RECT 71.785 18.075 71.955 18.245 ;
        RECT 71.785 12.635 71.955 12.805 ;
        RECT 72.245 56.155 72.415 56.325 ;
        RECT 72.245 50.715 72.415 50.885 ;
        RECT 72.245 45.275 72.415 45.445 ;
        RECT 72.245 39.835 72.415 40.005 ;
        RECT 72.245 34.395 72.415 34.565 ;
        RECT 72.245 28.955 72.415 29.125 ;
        RECT 72.245 23.515 72.415 23.685 ;
        RECT 72.245 18.075 72.415 18.245 ;
        RECT 72.245 12.635 72.415 12.805 ;
        RECT 72.705 56.155 72.875 56.325 ;
        RECT 72.705 50.715 72.875 50.885 ;
        RECT 72.705 45.275 72.875 45.445 ;
        RECT 72.705 39.835 72.875 40.005 ;
        RECT 72.705 34.395 72.875 34.565 ;
        RECT 72.705 28.955 72.875 29.125 ;
        RECT 72.705 23.515 72.875 23.685 ;
        RECT 72.705 18.075 72.875 18.245 ;
        RECT 72.705 12.635 72.875 12.805 ;
        RECT 73.165 56.155 73.335 56.325 ;
        RECT 73.165 50.715 73.335 50.885 ;
        RECT 73.165 45.275 73.335 45.445 ;
        RECT 73.165 39.835 73.335 40.005 ;
        RECT 73.165 34.395 73.335 34.565 ;
        RECT 73.165 28.955 73.335 29.125 ;
        RECT 73.165 23.515 73.335 23.685 ;
        RECT 73.165 18.075 73.335 18.245 ;
        RECT 73.165 12.635 73.335 12.805 ;
        RECT 73.625 56.155 73.795 56.325 ;
        RECT 73.625 50.715 73.795 50.885 ;
        RECT 73.625 45.275 73.795 45.445 ;
        RECT 73.625 39.835 73.795 40.005 ;
        RECT 73.625 34.395 73.795 34.565 ;
        RECT 73.625 28.955 73.795 29.125 ;
        RECT 73.625 23.515 73.795 23.685 ;
        RECT 73.625 18.075 73.795 18.245 ;
        RECT 73.625 12.635 73.795 12.805 ;
        RECT 74.085 56.155 74.255 56.325 ;
        RECT 74.085 50.715 74.255 50.885 ;
        RECT 74.085 45.275 74.255 45.445 ;
        RECT 74.085 39.835 74.255 40.005 ;
        RECT 74.085 34.395 74.255 34.565 ;
        RECT 74.085 28.955 74.255 29.125 ;
        RECT 74.085 23.515 74.255 23.685 ;
        RECT 74.085 18.075 74.255 18.245 ;
        RECT 74.085 12.635 74.255 12.805 ;
        RECT 74.545 56.155 74.715 56.325 ;
        RECT 74.545 50.715 74.715 50.885 ;
        RECT 74.545 45.275 74.715 45.445 ;
        RECT 74.545 39.835 74.715 40.005 ;
        RECT 74.545 34.395 74.715 34.565 ;
        RECT 74.545 28.955 74.715 29.125 ;
        RECT 74.545 23.515 74.715 23.685 ;
        RECT 74.545 18.075 74.715 18.245 ;
        RECT 74.545 12.635 74.715 12.805 ;
        RECT 75.005 56.155 75.175 56.325 ;
        RECT 75.005 50.715 75.175 50.885 ;
        RECT 75.005 45.275 75.175 45.445 ;
        RECT 75.005 39.835 75.175 40.005 ;
        RECT 75.005 34.395 75.175 34.565 ;
        RECT 75.005 28.955 75.175 29.125 ;
        RECT 75.005 23.515 75.175 23.685 ;
        RECT 75.005 18.075 75.175 18.245 ;
        RECT 75.005 12.635 75.175 12.805 ;
        RECT 75.465 56.155 75.635 56.325 ;
        RECT 75.465 50.715 75.635 50.885 ;
        RECT 75.465 45.275 75.635 45.445 ;
        RECT 75.465 39.835 75.635 40.005 ;
        RECT 75.465 34.395 75.635 34.565 ;
        RECT 75.465 28.955 75.635 29.125 ;
        RECT 75.465 23.515 75.635 23.685 ;
        RECT 75.465 18.075 75.635 18.245 ;
        RECT 75.465 12.635 75.635 12.805 ;
        RECT 75.925 56.155 76.095 56.325 ;
        RECT 75.925 50.715 76.095 50.885 ;
        RECT 75.925 45.275 76.095 45.445 ;
        RECT 75.925 39.835 76.095 40.005 ;
        RECT 75.925 34.395 76.095 34.565 ;
        RECT 75.925 28.955 76.095 29.125 ;
        RECT 75.925 23.515 76.095 23.685 ;
        RECT 75.925 18.075 76.095 18.245 ;
        RECT 75.925 12.635 76.095 12.805 ;
        RECT 76.385 56.155 76.555 56.325 ;
        RECT 76.385 50.715 76.555 50.885 ;
        RECT 76.385 45.275 76.555 45.445 ;
        RECT 76.385 39.835 76.555 40.005 ;
        RECT 76.385 34.395 76.555 34.565 ;
        RECT 76.385 28.955 76.555 29.125 ;
        RECT 76.385 23.515 76.555 23.685 ;
        RECT 76.385 18.075 76.555 18.245 ;
        RECT 76.385 12.635 76.555 12.805 ;
        RECT 76.845 56.155 77.015 56.325 ;
        RECT 76.845 50.715 77.015 50.885 ;
        RECT 76.845 45.275 77.015 45.445 ;
        RECT 76.845 39.835 77.015 40.005 ;
        RECT 76.845 34.395 77.015 34.565 ;
        RECT 76.845 28.955 77.015 29.125 ;
        RECT 76.845 23.515 77.015 23.685 ;
        RECT 76.845 18.075 77.015 18.245 ;
        RECT 76.845 12.635 77.015 12.805 ;
        RECT 77.305 56.155 77.475 56.325 ;
        RECT 77.305 50.715 77.475 50.885 ;
        RECT 77.305 45.275 77.475 45.445 ;
        RECT 77.305 39.835 77.475 40.005 ;
        RECT 77.305 34.395 77.475 34.565 ;
        RECT 77.305 28.955 77.475 29.125 ;
        RECT 77.305 23.515 77.475 23.685 ;
        RECT 77.305 18.075 77.475 18.245 ;
        RECT 77.305 12.635 77.475 12.805 ;
        RECT 77.765 56.155 77.935 56.325 ;
        RECT 77.765 50.715 77.935 50.885 ;
        RECT 77.765 45.275 77.935 45.445 ;
        RECT 77.765 39.835 77.935 40.005 ;
        RECT 77.765 34.395 77.935 34.565 ;
        RECT 77.765 28.955 77.935 29.125 ;
        RECT 77.765 23.515 77.935 23.685 ;
        RECT 77.765 18.075 77.935 18.245 ;
        RECT 77.765 12.635 77.935 12.805 ;
        RECT 78.225 56.155 78.395 56.325 ;
        RECT 78.225 50.715 78.395 50.885 ;
        RECT 78.225 45.275 78.395 45.445 ;
        RECT 78.225 39.835 78.395 40.005 ;
        RECT 78.225 34.395 78.395 34.565 ;
        RECT 78.225 28.955 78.395 29.125 ;
        RECT 78.225 23.515 78.395 23.685 ;
        RECT 78.225 18.075 78.395 18.245 ;
        RECT 78.225 12.635 78.395 12.805 ;
        RECT 78.685 56.155 78.855 56.325 ;
        RECT 78.685 50.715 78.855 50.885 ;
        RECT 78.685 45.275 78.855 45.445 ;
        RECT 78.685 39.835 78.855 40.005 ;
        RECT 78.685 34.395 78.855 34.565 ;
        RECT 78.685 28.955 78.855 29.125 ;
        RECT 78.685 23.515 78.855 23.685 ;
        RECT 78.685 18.075 78.855 18.245 ;
        RECT 78.685 12.635 78.855 12.805 ;
        RECT 79.145 56.155 79.315 56.325 ;
        RECT 79.145 50.715 79.315 50.885 ;
        RECT 79.145 45.275 79.315 45.445 ;
        RECT 79.145 39.835 79.315 40.005 ;
        RECT 79.145 34.395 79.315 34.565 ;
        RECT 79.145 28.955 79.315 29.125 ;
        RECT 79.145 23.515 79.315 23.685 ;
        RECT 79.145 18.075 79.315 18.245 ;
        RECT 79.145 12.635 79.315 12.805 ;
        RECT 79.605 56.155 79.775 56.325 ;
        RECT 79.605 50.715 79.775 50.885 ;
        RECT 79.605 45.275 79.775 45.445 ;
        RECT 79.605 39.835 79.775 40.005 ;
        RECT 79.605 34.395 79.775 34.565 ;
        RECT 79.605 28.955 79.775 29.125 ;
        RECT 79.605 23.515 79.775 23.685 ;
        RECT 79.605 18.075 79.775 18.245 ;
        RECT 79.605 12.635 79.775 12.805 ;
        RECT 80.065 56.155 80.235 56.325 ;
        RECT 80.065 50.715 80.235 50.885 ;
        RECT 80.065 45.275 80.235 45.445 ;
        RECT 80.065 39.835 80.235 40.005 ;
        RECT 80.065 34.395 80.235 34.565 ;
        RECT 80.065 28.955 80.235 29.125 ;
        RECT 80.065 23.515 80.235 23.685 ;
        RECT 80.065 18.075 80.235 18.245 ;
        RECT 80.065 12.635 80.235 12.805 ;
        RECT 80.525 56.155 80.695 56.325 ;
        RECT 80.525 50.715 80.695 50.885 ;
        RECT 80.525 45.275 80.695 45.445 ;
        RECT 80.525 39.835 80.695 40.005 ;
        RECT 80.525 34.395 80.695 34.565 ;
        RECT 80.525 28.955 80.695 29.125 ;
        RECT 80.525 23.515 80.695 23.685 ;
        RECT 80.525 18.075 80.695 18.245 ;
        RECT 80.525 12.635 80.695 12.805 ;
        RECT 80.985 56.155 81.155 56.325 ;
        RECT 80.985 50.715 81.155 50.885 ;
        RECT 80.985 45.275 81.155 45.445 ;
        RECT 80.985 39.835 81.155 40.005 ;
        RECT 80.985 34.395 81.155 34.565 ;
        RECT 80.985 28.955 81.155 29.125 ;
        RECT 80.985 23.515 81.155 23.685 ;
        RECT 80.985 18.075 81.155 18.245 ;
        RECT 80.985 12.635 81.155 12.805 ;
        RECT 81.445 56.155 81.615 56.325 ;
        RECT 81.445 50.715 81.615 50.885 ;
        RECT 81.445 45.275 81.615 45.445 ;
        RECT 81.445 39.835 81.615 40.005 ;
        RECT 81.445 34.395 81.615 34.565 ;
        RECT 81.445 28.955 81.615 29.125 ;
        RECT 81.445 23.515 81.615 23.685 ;
        RECT 81.445 18.075 81.615 18.245 ;
        RECT 81.445 12.635 81.615 12.805 ;
        RECT 81.905 56.155 82.075 56.325 ;
        RECT 81.905 50.715 82.075 50.885 ;
        RECT 81.905 45.275 82.075 45.445 ;
        RECT 81.905 39.835 82.075 40.005 ;
        RECT 81.905 34.395 82.075 34.565 ;
        RECT 81.905 28.955 82.075 29.125 ;
        RECT 81.905 23.515 82.075 23.685 ;
        RECT 81.905 18.075 82.075 18.245 ;
        RECT 81.905 12.635 82.075 12.805 ;
        RECT 82.365 56.155 82.535 56.325 ;
        RECT 82.365 50.715 82.535 50.885 ;
        RECT 82.365 45.275 82.535 45.445 ;
        RECT 82.365 39.835 82.535 40.005 ;
        RECT 82.365 34.395 82.535 34.565 ;
        RECT 82.365 28.955 82.535 29.125 ;
        RECT 82.365 23.515 82.535 23.685 ;
        RECT 82.365 18.075 82.535 18.245 ;
        RECT 82.365 12.635 82.535 12.805 ;
        RECT 82.825 56.155 82.995 56.325 ;
        RECT 82.825 50.715 82.995 50.885 ;
        RECT 82.825 45.275 82.995 45.445 ;
        RECT 82.825 39.835 82.995 40.005 ;
        RECT 82.825 34.395 82.995 34.565 ;
        RECT 82.825 28.955 82.995 29.125 ;
        RECT 82.825 23.515 82.995 23.685 ;
        RECT 82.825 18.075 82.995 18.245 ;
        RECT 82.825 12.635 82.995 12.805 ;
        RECT 83.285 56.155 83.455 56.325 ;
        RECT 83.285 50.715 83.455 50.885 ;
        RECT 83.285 45.275 83.455 45.445 ;
        RECT 83.285 39.835 83.455 40.005 ;
        RECT 83.285 34.395 83.455 34.565 ;
        RECT 83.285 28.955 83.455 29.125 ;
        RECT 83.285 23.515 83.455 23.685 ;
        RECT 83.285 18.075 83.455 18.245 ;
        RECT 83.285 12.635 83.455 12.805 ;
        RECT 83.745 56.155 83.915 56.325 ;
        RECT 83.745 50.715 83.915 50.885 ;
        RECT 83.745 45.275 83.915 45.445 ;
        RECT 83.745 39.835 83.915 40.005 ;
        RECT 83.745 34.395 83.915 34.565 ;
        RECT 83.745 28.955 83.915 29.125 ;
        RECT 83.745 23.515 83.915 23.685 ;
        RECT 83.745 18.075 83.915 18.245 ;
        RECT 83.745 12.635 83.915 12.805 ;
        RECT 84.205 56.155 84.375 56.325 ;
        RECT 84.205 50.715 84.375 50.885 ;
        RECT 84.205 45.275 84.375 45.445 ;
        RECT 84.205 39.835 84.375 40.005 ;
        RECT 84.205 34.395 84.375 34.565 ;
        RECT 84.205 28.955 84.375 29.125 ;
        RECT 84.205 23.515 84.375 23.685 ;
        RECT 84.205 18.075 84.375 18.245 ;
        RECT 84.205 12.635 84.375 12.805 ;
        RECT 84.665 56.155 84.835 56.325 ;
        RECT 84.665 50.715 84.835 50.885 ;
        RECT 84.665 45.275 84.835 45.445 ;
        RECT 84.665 39.835 84.835 40.005 ;
        RECT 84.665 34.395 84.835 34.565 ;
        RECT 84.665 28.955 84.835 29.125 ;
        RECT 84.665 23.515 84.835 23.685 ;
        RECT 84.665 18.075 84.835 18.245 ;
        RECT 84.665 12.635 84.835 12.805 ;
        RECT 85.125 56.155 85.295 56.325 ;
        RECT 85.125 50.715 85.295 50.885 ;
        RECT 85.125 45.275 85.295 45.445 ;
        RECT 85.125 39.835 85.295 40.005 ;
        RECT 85.125 34.395 85.295 34.565 ;
        RECT 85.125 28.955 85.295 29.125 ;
        RECT 85.125 23.515 85.295 23.685 ;
        RECT 85.125 18.075 85.295 18.245 ;
        RECT 85.125 12.635 85.295 12.805 ;
        RECT 85.585 56.155 85.755 56.325 ;
        RECT 85.585 50.715 85.755 50.885 ;
        RECT 85.585 45.275 85.755 45.445 ;
        RECT 85.585 39.835 85.755 40.005 ;
        RECT 85.585 34.395 85.755 34.565 ;
        RECT 85.585 28.955 85.755 29.125 ;
        RECT 85.585 23.515 85.755 23.685 ;
        RECT 85.585 18.075 85.755 18.245 ;
        RECT 85.585 12.635 85.755 12.805 ;
        RECT 86.045 56.155 86.215 56.325 ;
        RECT 86.045 50.715 86.215 50.885 ;
        RECT 86.045 45.275 86.215 45.445 ;
        RECT 86.045 39.835 86.215 40.005 ;
        RECT 86.045 34.395 86.215 34.565 ;
        RECT 86.045 28.955 86.215 29.125 ;
        RECT 86.045 23.515 86.215 23.685 ;
        RECT 86.045 18.075 86.215 18.245 ;
        RECT 86.045 12.635 86.215 12.805 ;
        RECT 86.505 56.155 86.675 56.325 ;
        RECT 86.505 50.715 86.675 50.885 ;
        RECT 86.505 45.275 86.675 45.445 ;
        RECT 86.505 39.835 86.675 40.005 ;
        RECT 86.505 34.395 86.675 34.565 ;
        RECT 86.505 28.955 86.675 29.125 ;
        RECT 86.505 23.515 86.675 23.685 ;
        RECT 86.505 18.075 86.675 18.245 ;
        RECT 86.505 12.635 86.675 12.805 ;
        RECT 86.965 56.155 87.135 56.325 ;
        RECT 86.965 50.715 87.135 50.885 ;
        RECT 86.965 45.275 87.135 45.445 ;
        RECT 86.965 39.835 87.135 40.005 ;
        RECT 86.965 34.395 87.135 34.565 ;
        RECT 86.965 28.955 87.135 29.125 ;
        RECT 86.965 23.515 87.135 23.685 ;
        RECT 86.965 18.075 87.135 18.245 ;
        RECT 86.965 12.635 87.135 12.805 ;
        RECT 87.425 56.155 87.595 56.325 ;
        RECT 87.425 50.715 87.595 50.885 ;
        RECT 87.425 45.275 87.595 45.445 ;
        RECT 87.425 39.835 87.595 40.005 ;
        RECT 87.425 34.395 87.595 34.565 ;
        RECT 87.425 28.955 87.595 29.125 ;
        RECT 87.425 23.515 87.595 23.685 ;
        RECT 87.425 18.075 87.595 18.245 ;
        RECT 87.425 12.635 87.595 12.805 ;
        RECT 87.885 56.155 88.055 56.325 ;
        RECT 87.885 50.715 88.055 50.885 ;
        RECT 87.885 45.275 88.055 45.445 ;
        RECT 87.885 39.835 88.055 40.005 ;
        RECT 87.885 34.395 88.055 34.565 ;
        RECT 87.885 28.955 88.055 29.125 ;
        RECT 87.885 23.515 88.055 23.685 ;
        RECT 87.885 18.075 88.055 18.245 ;
        RECT 87.885 12.635 88.055 12.805 ;
        RECT 88.345 56.155 88.515 56.325 ;
        RECT 88.345 50.715 88.515 50.885 ;
        RECT 88.345 45.275 88.515 45.445 ;
        RECT 88.345 39.835 88.515 40.005 ;
        RECT 88.345 34.395 88.515 34.565 ;
        RECT 88.345 28.955 88.515 29.125 ;
        RECT 88.345 23.515 88.515 23.685 ;
        RECT 88.345 18.075 88.515 18.245 ;
        RECT 88.345 12.635 88.515 12.805 ;
        RECT 88.805 56.155 88.975 56.325 ;
        RECT 88.805 50.715 88.975 50.885 ;
        RECT 88.805 45.275 88.975 45.445 ;
        RECT 88.805 39.835 88.975 40.005 ;
        RECT 88.805 34.395 88.975 34.565 ;
        RECT 88.805 28.955 88.975 29.125 ;
        RECT 88.805 23.515 88.975 23.685 ;
        RECT 88.805 18.075 88.975 18.245 ;
        RECT 88.805 12.635 88.975 12.805 ;
        RECT 89.265 56.155 89.435 56.325 ;
        RECT 89.265 50.715 89.435 50.885 ;
        RECT 89.265 45.275 89.435 45.445 ;
        RECT 89.265 39.835 89.435 40.005 ;
        RECT 89.265 34.395 89.435 34.565 ;
        RECT 89.265 28.955 89.435 29.125 ;
        RECT 89.265 23.515 89.435 23.685 ;
        RECT 89.265 18.075 89.435 18.245 ;
        RECT 89.265 12.635 89.435 12.805 ;
        RECT 89.725 56.155 89.895 56.325 ;
        RECT 89.725 50.715 89.895 50.885 ;
        RECT 89.725 45.275 89.895 45.445 ;
        RECT 89.725 39.835 89.895 40.005 ;
        RECT 89.725 34.395 89.895 34.565 ;
        RECT 89.725 28.955 89.895 29.125 ;
        RECT 89.725 23.515 89.895 23.685 ;
        RECT 89.725 18.075 89.895 18.245 ;
        RECT 89.725 12.635 89.895 12.805 ;
        RECT 90.185 56.155 90.355 56.325 ;
        RECT 90.185 50.715 90.355 50.885 ;
        RECT 90.185 45.275 90.355 45.445 ;
        RECT 90.185 39.835 90.355 40.005 ;
        RECT 90.185 34.395 90.355 34.565 ;
        RECT 90.185 28.955 90.355 29.125 ;
        RECT 90.185 23.515 90.355 23.685 ;
        RECT 90.185 18.075 90.355 18.245 ;
        RECT 90.185 12.635 90.355 12.805 ;
        RECT 90.645 56.155 90.815 56.325 ;
        RECT 90.645 50.715 90.815 50.885 ;
        RECT 90.645 45.275 90.815 45.445 ;
        RECT 90.645 39.835 90.815 40.005 ;
        RECT 90.645 34.395 90.815 34.565 ;
        RECT 90.645 28.955 90.815 29.125 ;
        RECT 90.645 23.515 90.815 23.685 ;
        RECT 90.645 18.075 90.815 18.245 ;
        RECT 90.645 12.635 90.815 12.805 ;
        RECT 91.105 56.155 91.275 56.325 ;
        RECT 91.105 50.715 91.275 50.885 ;
        RECT 91.105 45.275 91.275 45.445 ;
        RECT 91.105 39.835 91.275 40.005 ;
        RECT 91.105 34.395 91.275 34.565 ;
        RECT 91.105 28.955 91.275 29.125 ;
        RECT 91.105 23.515 91.275 23.685 ;
        RECT 91.105 18.075 91.275 18.245 ;
        RECT 91.105 12.635 91.275 12.805 ;
        RECT 91.565 56.155 91.735 56.325 ;
        RECT 91.565 50.715 91.735 50.885 ;
        RECT 91.565 45.275 91.735 45.445 ;
        RECT 91.565 39.835 91.735 40.005 ;
        RECT 91.565 34.395 91.735 34.565 ;
        RECT 91.565 28.955 91.735 29.125 ;
        RECT 91.565 23.515 91.735 23.685 ;
        RECT 91.565 18.075 91.735 18.245 ;
        RECT 91.565 12.635 91.735 12.805 ;
        RECT 92.025 56.155 92.195 56.325 ;
        RECT 92.025 50.715 92.195 50.885 ;
        RECT 92.025 45.275 92.195 45.445 ;
        RECT 92.025 39.835 92.195 40.005 ;
        RECT 92.025 34.395 92.195 34.565 ;
        RECT 92.025 28.955 92.195 29.125 ;
        RECT 92.025 23.515 92.195 23.685 ;
        RECT 92.025 18.075 92.195 18.245 ;
        RECT 92.025 12.635 92.195 12.805 ;
        RECT 92.485 56.155 92.655 56.325 ;
        RECT 92.485 50.715 92.655 50.885 ;
        RECT 92.485 45.275 92.655 45.445 ;
        RECT 92.485 39.835 92.655 40.005 ;
        RECT 92.485 34.395 92.655 34.565 ;
        RECT 92.485 28.955 92.655 29.125 ;
        RECT 92.485 23.515 92.655 23.685 ;
        RECT 92.485 18.075 92.655 18.245 ;
        RECT 92.485 12.635 92.655 12.805 ;
        RECT 92.945 56.155 93.115 56.325 ;
        RECT 92.945 50.715 93.115 50.885 ;
        RECT 92.945 45.275 93.115 45.445 ;
        RECT 92.945 39.835 93.115 40.005 ;
        RECT 92.945 34.395 93.115 34.565 ;
        RECT 92.945 28.955 93.115 29.125 ;
        RECT 92.945 23.515 93.115 23.685 ;
        RECT 92.945 18.075 93.115 18.245 ;
        RECT 92.945 12.635 93.115 12.805 ;
        RECT 93.405 56.155 93.575 56.325 ;
        RECT 93.405 50.715 93.575 50.885 ;
        RECT 93.405 45.275 93.575 45.445 ;
        RECT 93.405 39.835 93.575 40.005 ;
        RECT 93.405 34.395 93.575 34.565 ;
        RECT 93.405 28.955 93.575 29.125 ;
        RECT 93.405 23.515 93.575 23.685 ;
        RECT 93.405 18.075 93.575 18.245 ;
        RECT 93.405 12.635 93.575 12.805 ;
        RECT 93.865 56.155 94.035 56.325 ;
        RECT 93.865 50.715 94.035 50.885 ;
        RECT 93.865 45.275 94.035 45.445 ;
        RECT 93.865 39.835 94.035 40.005 ;
        RECT 93.865 34.395 94.035 34.565 ;
        RECT 93.865 28.955 94.035 29.125 ;
        RECT 93.865 23.515 94.035 23.685 ;
        RECT 93.865 18.075 94.035 18.245 ;
        RECT 93.865 12.635 94.035 12.805 ;
        RECT 94.325 56.155 94.495 56.325 ;
        RECT 94.325 50.715 94.495 50.885 ;
        RECT 94.325 45.275 94.495 45.445 ;
        RECT 94.325 39.835 94.495 40.005 ;
        RECT 94.325 34.395 94.495 34.565 ;
        RECT 94.325 28.955 94.495 29.125 ;
        RECT 94.325 23.515 94.495 23.685 ;
        RECT 94.325 18.075 94.495 18.245 ;
        RECT 94.325 12.635 94.495 12.805 ;
        RECT 94.785 56.155 94.955 56.325 ;
        RECT 94.785 50.715 94.955 50.885 ;
        RECT 94.785 45.275 94.955 45.445 ;
        RECT 94.785 39.835 94.955 40.005 ;
        RECT 94.785 34.395 94.955 34.565 ;
        RECT 94.785 28.955 94.955 29.125 ;
        RECT 94.785 23.515 94.955 23.685 ;
        RECT 94.785 18.075 94.955 18.245 ;
        RECT 94.785 12.635 94.955 12.805 ;
        RECT 95.245 56.155 95.415 56.325 ;
        RECT 95.245 50.715 95.415 50.885 ;
        RECT 95.245 45.275 95.415 45.445 ;
        RECT 95.245 39.835 95.415 40.005 ;
        RECT 95.245 34.395 95.415 34.565 ;
        RECT 95.245 28.955 95.415 29.125 ;
        RECT 95.245 23.515 95.415 23.685 ;
        RECT 95.245 18.075 95.415 18.245 ;
        RECT 95.245 12.635 95.415 12.805 ;
        RECT 95.705 56.155 95.875 56.325 ;
        RECT 95.705 50.715 95.875 50.885 ;
        RECT 95.705 45.275 95.875 45.445 ;
        RECT 95.705 39.835 95.875 40.005 ;
        RECT 95.705 34.395 95.875 34.565 ;
        RECT 95.705 28.955 95.875 29.125 ;
        RECT 95.705 23.515 95.875 23.685 ;
        RECT 95.705 18.075 95.875 18.245 ;
        RECT 95.705 12.635 95.875 12.805 ;
        RECT 96.165 56.155 96.335 56.325 ;
        RECT 96.165 50.715 96.335 50.885 ;
        RECT 96.165 45.275 96.335 45.445 ;
        RECT 96.165 39.835 96.335 40.005 ;
        RECT 96.165 34.395 96.335 34.565 ;
        RECT 96.165 28.955 96.335 29.125 ;
        RECT 96.165 23.515 96.335 23.685 ;
        RECT 96.165 18.075 96.335 18.245 ;
        RECT 96.165 12.635 96.335 12.805 ;
        RECT 96.625 56.155 96.795 56.325 ;
        RECT 96.625 50.715 96.795 50.885 ;
        RECT 96.625 45.275 96.795 45.445 ;
        RECT 96.625 39.835 96.795 40.005 ;
        RECT 96.625 34.395 96.795 34.565 ;
        RECT 96.625 28.955 96.795 29.125 ;
        RECT 96.625 23.515 96.795 23.685 ;
        RECT 96.625 18.075 96.795 18.245 ;
        RECT 96.625 12.635 96.795 12.805 ;
        RECT 97.085 56.155 97.255 56.325 ;
        RECT 97.085 50.715 97.255 50.885 ;
        RECT 97.085 45.275 97.255 45.445 ;
        RECT 97.085 39.835 97.255 40.005 ;
        RECT 97.085 34.395 97.255 34.565 ;
        RECT 97.085 28.955 97.255 29.125 ;
        RECT 97.085 23.515 97.255 23.685 ;
        RECT 97.085 18.075 97.255 18.245 ;
        RECT 97.085 12.635 97.255 12.805 ;
        RECT 97.545 56.155 97.715 56.325 ;
        RECT 97.545 50.715 97.715 50.885 ;
        RECT 97.545 45.275 97.715 45.445 ;
        RECT 97.545 39.835 97.715 40.005 ;
        RECT 97.545 34.395 97.715 34.565 ;
        RECT 97.545 28.955 97.715 29.125 ;
        RECT 97.545 23.515 97.715 23.685 ;
        RECT 97.545 18.075 97.715 18.245 ;
        RECT 97.545 12.635 97.715 12.805 ;
        RECT 98.005 56.155 98.175 56.325 ;
        RECT 98.005 50.715 98.175 50.885 ;
        RECT 98.005 45.275 98.175 45.445 ;
        RECT 98.005 39.835 98.175 40.005 ;
        RECT 98.005 34.395 98.175 34.565 ;
        RECT 98.005 28.955 98.175 29.125 ;
        RECT 98.005 23.515 98.175 23.685 ;
        RECT 98.005 18.075 98.175 18.245 ;
        RECT 98.005 12.635 98.175 12.805 ;
        RECT 98.465 56.155 98.635 56.325 ;
        RECT 98.465 50.715 98.635 50.885 ;
        RECT 98.465 45.275 98.635 45.445 ;
        RECT 98.465 39.835 98.635 40.005 ;
        RECT 98.465 34.395 98.635 34.565 ;
        RECT 98.465 28.955 98.635 29.125 ;
        RECT 98.465 23.515 98.635 23.685 ;
        RECT 98.465 18.075 98.635 18.245 ;
        RECT 98.465 12.635 98.635 12.805 ;
        RECT 98.925 56.155 99.095 56.325 ;
        RECT 98.925 50.715 99.095 50.885 ;
        RECT 98.925 45.275 99.095 45.445 ;
        RECT 98.925 39.835 99.095 40.005 ;
        RECT 98.925 34.395 99.095 34.565 ;
        RECT 98.925 28.955 99.095 29.125 ;
        RECT 98.925 23.515 99.095 23.685 ;
        RECT 98.925 18.075 99.095 18.245 ;
        RECT 98.925 12.635 99.095 12.805 ;
        RECT 99.385 56.155 99.555 56.325 ;
        RECT 99.385 50.715 99.555 50.885 ;
        RECT 99.385 45.275 99.555 45.445 ;
        RECT 99.385 39.835 99.555 40.005 ;
        RECT 99.385 34.395 99.555 34.565 ;
        RECT 99.385 28.955 99.555 29.125 ;
        RECT 99.385 23.515 99.555 23.685 ;
        RECT 99.385 18.075 99.555 18.245 ;
        RECT 99.385 12.635 99.555 12.805 ;
        RECT 99.845 56.155 100.015 56.325 ;
        RECT 99.845 50.715 100.015 50.885 ;
        RECT 99.845 45.275 100.015 45.445 ;
        RECT 99.845 39.835 100.015 40.005 ;
        RECT 99.845 34.395 100.015 34.565 ;
        RECT 99.845 28.955 100.015 29.125 ;
        RECT 99.845 23.515 100.015 23.685 ;
        RECT 99.845 18.075 100.015 18.245 ;
        RECT 99.845 12.635 100.015 12.805 ;
        RECT 100.305 56.155 100.475 56.325 ;
        RECT 100.305 50.715 100.475 50.885 ;
        RECT 100.305 45.275 100.475 45.445 ;
        RECT 100.305 39.835 100.475 40.005 ;
        RECT 100.305 34.395 100.475 34.565 ;
        RECT 100.305 28.955 100.475 29.125 ;
        RECT 100.305 23.515 100.475 23.685 ;
        RECT 100.305 18.075 100.475 18.245 ;
        RECT 100.305 12.635 100.475 12.805 ;
        RECT 100.765 56.155 100.935 56.325 ;
        RECT 100.765 50.715 100.935 50.885 ;
        RECT 100.765 45.275 100.935 45.445 ;
        RECT 100.765 39.835 100.935 40.005 ;
        RECT 100.765 34.395 100.935 34.565 ;
        RECT 100.765 28.955 100.935 29.125 ;
        RECT 100.765 23.515 100.935 23.685 ;
        RECT 100.765 18.075 100.935 18.245 ;
        RECT 100.765 12.635 100.935 12.805 ;
        RECT 101.225 56.155 101.395 56.325 ;
        RECT 101.225 50.715 101.395 50.885 ;
        RECT 101.225 45.275 101.395 45.445 ;
        RECT 101.225 39.835 101.395 40.005 ;
        RECT 101.225 34.395 101.395 34.565 ;
        RECT 101.225 28.955 101.395 29.125 ;
        RECT 101.225 23.515 101.395 23.685 ;
        RECT 101.225 18.075 101.395 18.245 ;
        RECT 101.225 12.635 101.395 12.805 ;
        RECT 101.685 56.155 101.855 56.325 ;
        RECT 101.685 50.715 101.855 50.885 ;
        RECT 101.685 45.275 101.855 45.445 ;
        RECT 101.685 39.835 101.855 40.005 ;
        RECT 101.685 34.395 101.855 34.565 ;
        RECT 101.685 28.955 101.855 29.125 ;
        RECT 101.685 23.515 101.855 23.685 ;
        RECT 101.685 18.075 101.855 18.245 ;
        RECT 101.685 12.635 101.855 12.805 ;
        RECT 102.145 56.155 102.315 56.325 ;
        RECT 102.145 50.715 102.315 50.885 ;
        RECT 102.145 45.275 102.315 45.445 ;
        RECT 102.145 39.835 102.315 40.005 ;
        RECT 102.145 34.395 102.315 34.565 ;
        RECT 102.145 28.955 102.315 29.125 ;
        RECT 102.145 23.515 102.315 23.685 ;
        RECT 102.145 18.075 102.315 18.245 ;
        RECT 102.145 12.635 102.315 12.805 ;
        RECT 102.605 56.155 102.775 56.325 ;
        RECT 102.605 50.715 102.775 50.885 ;
        RECT 102.605 45.275 102.775 45.445 ;
        RECT 102.605 39.835 102.775 40.005 ;
        RECT 102.605 34.395 102.775 34.565 ;
        RECT 102.605 28.955 102.775 29.125 ;
        RECT 102.605 23.515 102.775 23.685 ;
        RECT 102.605 18.075 102.775 18.245 ;
        RECT 102.605 12.635 102.775 12.805 ;
        RECT 103.065 56.155 103.235 56.325 ;
        RECT 103.065 50.715 103.235 50.885 ;
        RECT 103.065 45.275 103.235 45.445 ;
        RECT 103.065 39.835 103.235 40.005 ;
        RECT 103.065 34.395 103.235 34.565 ;
        RECT 103.065 28.955 103.235 29.125 ;
        RECT 103.065 23.515 103.235 23.685 ;
        RECT 103.065 18.075 103.235 18.245 ;
        RECT 103.065 12.635 103.235 12.805 ;
        RECT 103.525 56.155 103.695 56.325 ;
        RECT 103.525 50.715 103.695 50.885 ;
        RECT 103.525 45.275 103.695 45.445 ;
        RECT 103.525 39.835 103.695 40.005 ;
        RECT 103.525 34.395 103.695 34.565 ;
        RECT 103.525 28.955 103.695 29.125 ;
        RECT 103.525 23.515 103.695 23.685 ;
        RECT 103.525 18.075 103.695 18.245 ;
        RECT 103.525 12.635 103.695 12.805 ;
        RECT 103.985 56.155 104.155 56.325 ;
        RECT 103.985 50.715 104.155 50.885 ;
        RECT 103.985 45.275 104.155 45.445 ;
        RECT 103.985 39.835 104.155 40.005 ;
        RECT 103.985 34.395 104.155 34.565 ;
        RECT 103.985 28.955 104.155 29.125 ;
        RECT 103.985 23.515 104.155 23.685 ;
        RECT 103.985 18.075 104.155 18.245 ;
        RECT 103.985 12.635 104.155 12.805 ;
        RECT 104.445 56.155 104.615 56.325 ;
        RECT 104.445 50.715 104.615 50.885 ;
        RECT 104.445 45.275 104.615 45.445 ;
        RECT 104.445 39.835 104.615 40.005 ;
        RECT 104.445 34.395 104.615 34.565 ;
        RECT 104.445 28.955 104.615 29.125 ;
        RECT 104.445 23.515 104.615 23.685 ;
        RECT 104.445 18.075 104.615 18.245 ;
        RECT 104.445 12.635 104.615 12.805 ;
        RECT 104.905 56.155 105.075 56.325 ;
        RECT 104.905 50.715 105.075 50.885 ;
        RECT 104.905 45.275 105.075 45.445 ;
        RECT 104.905 39.835 105.075 40.005 ;
        RECT 104.905 34.395 105.075 34.565 ;
        RECT 104.905 28.955 105.075 29.125 ;
        RECT 104.905 23.515 105.075 23.685 ;
        RECT 104.905 18.075 105.075 18.245 ;
        RECT 104.905 12.635 105.075 12.805 ;
        RECT 105.365 56.155 105.535 56.325 ;
        RECT 105.365 50.715 105.535 50.885 ;
        RECT 105.365 45.275 105.535 45.445 ;
        RECT 105.365 39.835 105.535 40.005 ;
        RECT 105.365 34.395 105.535 34.565 ;
        RECT 105.365 28.955 105.535 29.125 ;
        RECT 105.365 23.515 105.535 23.685 ;
        RECT 105.365 18.075 105.535 18.245 ;
        RECT 105.365 12.635 105.535 12.805 ;
        RECT 105.825 56.155 105.995 56.325 ;
        RECT 105.825 50.715 105.995 50.885 ;
        RECT 105.825 45.275 105.995 45.445 ;
        RECT 105.825 39.835 105.995 40.005 ;
        RECT 105.825 34.395 105.995 34.565 ;
        RECT 105.825 28.955 105.995 29.125 ;
        RECT 105.825 23.515 105.995 23.685 ;
        RECT 105.825 18.075 105.995 18.245 ;
        RECT 105.825 12.635 105.995 12.805 ;
        RECT 106.285 56.155 106.455 56.325 ;
        RECT 106.285 50.715 106.455 50.885 ;
        RECT 106.285 45.275 106.455 45.445 ;
        RECT 106.285 39.835 106.455 40.005 ;
        RECT 106.285 34.395 106.455 34.565 ;
        RECT 106.285 28.955 106.455 29.125 ;
        RECT 106.285 23.515 106.455 23.685 ;
        RECT 106.285 18.075 106.455 18.245 ;
        RECT 106.285 12.635 106.455 12.805 ;
        RECT 106.745 56.155 106.915 56.325 ;
        RECT 106.745 50.715 106.915 50.885 ;
        RECT 106.745 45.275 106.915 45.445 ;
        RECT 106.745 39.835 106.915 40.005 ;
        RECT 106.745 34.395 106.915 34.565 ;
        RECT 106.745 28.955 106.915 29.125 ;
        RECT 106.745 23.515 106.915 23.685 ;
        RECT 106.745 18.075 106.915 18.245 ;
        RECT 106.745 12.635 106.915 12.805 ;
        RECT 107.205 56.155 107.375 56.325 ;
        RECT 107.205 50.715 107.375 50.885 ;
        RECT 107.205 45.275 107.375 45.445 ;
        RECT 107.205 39.835 107.375 40.005 ;
        RECT 107.205 34.395 107.375 34.565 ;
        RECT 107.205 28.955 107.375 29.125 ;
        RECT 107.205 23.515 107.375 23.685 ;
        RECT 107.205 18.075 107.375 18.245 ;
        RECT 107.205 12.635 107.375 12.805 ;
        RECT 107.665 56.155 107.835 56.325 ;
        RECT 107.665 50.715 107.835 50.885 ;
        RECT 107.665 45.275 107.835 45.445 ;
        RECT 107.665 39.835 107.835 40.005 ;
        RECT 107.665 34.395 107.835 34.565 ;
        RECT 107.665 28.955 107.835 29.125 ;
        RECT 107.665 23.515 107.835 23.685 ;
        RECT 107.665 18.075 107.835 18.245 ;
        RECT 107.665 12.635 107.835 12.805 ;
        RECT 108.125 56.155 108.295 56.325 ;
        RECT 108.125 50.715 108.295 50.885 ;
        RECT 108.125 45.275 108.295 45.445 ;
        RECT 108.125 39.835 108.295 40.005 ;
        RECT 108.125 34.395 108.295 34.565 ;
        RECT 108.125 28.955 108.295 29.125 ;
        RECT 108.125 23.515 108.295 23.685 ;
        RECT 108.125 18.075 108.295 18.245 ;
        RECT 108.125 12.635 108.295 12.805 ;
        RECT 108.585 56.155 108.755 56.325 ;
        RECT 108.585 50.715 108.755 50.885 ;
        RECT 108.585 45.275 108.755 45.445 ;
        RECT 108.585 39.835 108.755 40.005 ;
        RECT 108.585 34.395 108.755 34.565 ;
        RECT 108.585 28.955 108.755 29.125 ;
        RECT 108.585 23.515 108.755 23.685 ;
        RECT 108.585 18.075 108.755 18.245 ;
        RECT 108.585 12.635 108.755 12.805 ;
        RECT 109.045 56.155 109.215 56.325 ;
        RECT 109.045 50.715 109.215 50.885 ;
        RECT 109.045 45.275 109.215 45.445 ;
        RECT 109.045 39.835 109.215 40.005 ;
        RECT 109.045 34.395 109.215 34.565 ;
        RECT 109.045 28.955 109.215 29.125 ;
        RECT 109.045 23.515 109.215 23.685 ;
        RECT 109.045 18.075 109.215 18.245 ;
        RECT 109.045 12.635 109.215 12.805 ;
        RECT 109.505 56.155 109.675 56.325 ;
        RECT 109.505 50.715 109.675 50.885 ;
        RECT 109.505 45.275 109.675 45.445 ;
        RECT 109.505 39.835 109.675 40.005 ;
        RECT 109.505 34.395 109.675 34.565 ;
        RECT 109.505 28.955 109.675 29.125 ;
        RECT 109.505 23.515 109.675 23.685 ;
        RECT 109.505 18.075 109.675 18.245 ;
        RECT 109.505 12.635 109.675 12.805 ;
        RECT 109.965 56.155 110.135 56.325 ;
        RECT 109.965 50.715 110.135 50.885 ;
        RECT 109.965 45.275 110.135 45.445 ;
        RECT 109.965 39.835 110.135 40.005 ;
        RECT 109.965 34.395 110.135 34.565 ;
        RECT 109.965 28.955 110.135 29.125 ;
        RECT 109.965 23.515 110.135 23.685 ;
        RECT 109.965 18.075 110.135 18.245 ;
        RECT 109.965 12.635 110.135 12.805 ;
        RECT 110.425 56.155 110.595 56.325 ;
        RECT 110.425 50.715 110.595 50.885 ;
        RECT 110.425 45.275 110.595 45.445 ;
        RECT 110.425 39.835 110.595 40.005 ;
        RECT 110.425 34.395 110.595 34.565 ;
        RECT 110.425 28.955 110.595 29.125 ;
        RECT 110.425 23.515 110.595 23.685 ;
        RECT 110.425 18.075 110.595 18.245 ;
        RECT 110.425 12.635 110.595 12.805 ;
        RECT 110.885 56.155 111.055 56.325 ;
        RECT 110.885 50.715 111.055 50.885 ;
        RECT 110.885 45.275 111.055 45.445 ;
        RECT 110.885 39.835 111.055 40.005 ;
        RECT 110.885 34.395 111.055 34.565 ;
        RECT 110.885 28.955 111.055 29.125 ;
        RECT 110.885 23.515 111.055 23.685 ;
        RECT 110.885 18.075 111.055 18.245 ;
        RECT 110.885 12.635 111.055 12.805 ;
        RECT 111.345 56.155 111.515 56.325 ;
        RECT 111.345 50.715 111.515 50.885 ;
        RECT 111.345 45.275 111.515 45.445 ;
        RECT 111.345 39.835 111.515 40.005 ;
        RECT 111.345 34.395 111.515 34.565 ;
        RECT 111.345 28.955 111.515 29.125 ;
        RECT 111.345 23.515 111.515 23.685 ;
        RECT 111.345 18.075 111.515 18.245 ;
        RECT 111.345 12.635 111.515 12.805 ;
        RECT 111.805 56.155 111.975 56.325 ;
        RECT 111.805 50.715 111.975 50.885 ;
        RECT 111.805 45.275 111.975 45.445 ;
        RECT 111.805 39.835 111.975 40.005 ;
        RECT 111.805 34.395 111.975 34.565 ;
        RECT 111.805 28.955 111.975 29.125 ;
        RECT 111.805 23.515 111.975 23.685 ;
        RECT 111.805 18.075 111.975 18.245 ;
        RECT 111.805 12.635 111.975 12.805 ;
        RECT 112.265 56.155 112.435 56.325 ;
        RECT 112.265 50.715 112.435 50.885 ;
        RECT 10.145 56.155 10.315 56.325 ;
        RECT 10.145 50.715 10.315 50.885 ;
        RECT 10.145 45.275 10.315 45.445 ;
        RECT 10.145 39.835 10.315 40.005 ;
        RECT 10.145 34.395 10.315 34.565 ;
        RECT 10.145 28.955 10.315 29.125 ;
        RECT 10.145 23.515 10.315 23.685 ;
        RECT 10.145 18.075 10.315 18.245 ;
        RECT 10.145 12.635 10.315 12.805 ;
        RECT 10.605 56.155 10.775 56.325 ;
        RECT 10.605 50.715 10.775 50.885 ;
        RECT 10.605 45.275 10.775 45.445 ;
        RECT 10.605 39.835 10.775 40.005 ;
        RECT 10.605 34.395 10.775 34.565 ;
        RECT 10.605 28.955 10.775 29.125 ;
        RECT 10.605 23.515 10.775 23.685 ;
        RECT 10.605 18.075 10.775 18.245 ;
        RECT 10.605 12.635 10.775 12.805 ;
        RECT 11.065 56.155 11.235 56.325 ;
        RECT 11.065 50.715 11.235 50.885 ;
        RECT 11.065 45.275 11.235 45.445 ;
        RECT 11.065 39.835 11.235 40.005 ;
        RECT 11.065 34.395 11.235 34.565 ;
        RECT 11.065 28.955 11.235 29.125 ;
        RECT 11.065 23.515 11.235 23.685 ;
        RECT 11.065 18.075 11.235 18.245 ;
        RECT 11.065 12.635 11.235 12.805 ;
        RECT 11.525 56.155 11.695 56.325 ;
        RECT 11.525 50.715 11.695 50.885 ;
        RECT 11.525 45.275 11.695 45.445 ;
        RECT 11.525 39.835 11.695 40.005 ;
        RECT 11.525 34.395 11.695 34.565 ;
        RECT 11.525 28.955 11.695 29.125 ;
        RECT 11.525 23.515 11.695 23.685 ;
        RECT 11.525 18.075 11.695 18.245 ;
        RECT 11.525 12.635 11.695 12.805 ;
        RECT 11.985 56.155 12.155 56.325 ;
        RECT 11.985 50.715 12.155 50.885 ;
        RECT 11.985 45.275 12.155 45.445 ;
        RECT 11.985 39.835 12.155 40.005 ;
        RECT 11.985 34.395 12.155 34.565 ;
        RECT 11.985 28.955 12.155 29.125 ;
        RECT 11.985 23.515 12.155 23.685 ;
        RECT 11.985 18.075 12.155 18.245 ;
        RECT 11.985 12.635 12.155 12.805 ;
        RECT 12.445 56.155 12.615 56.325 ;
        RECT 12.445 50.715 12.615 50.885 ;
        RECT 12.445 45.275 12.615 45.445 ;
        RECT 12.445 39.835 12.615 40.005 ;
        RECT 12.445 34.395 12.615 34.565 ;
        RECT 12.445 28.955 12.615 29.125 ;
        RECT 12.445 23.515 12.615 23.685 ;
        RECT 12.445 18.075 12.615 18.245 ;
        RECT 12.445 12.635 12.615 12.805 ;
        RECT 12.905 56.155 13.075 56.325 ;
        RECT 12.905 50.715 13.075 50.885 ;
        RECT 12.905 45.275 13.075 45.445 ;
        RECT 12.905 39.835 13.075 40.005 ;
        RECT 12.905 34.395 13.075 34.565 ;
        RECT 12.905 28.955 13.075 29.125 ;
        RECT 12.905 23.515 13.075 23.685 ;
        RECT 12.905 18.075 13.075 18.245 ;
        RECT 12.905 12.635 13.075 12.805 ;
        RECT 13.365 56.155 13.535 56.325 ;
        RECT 13.365 50.715 13.535 50.885 ;
        RECT 13.365 45.275 13.535 45.445 ;
        RECT 13.365 39.835 13.535 40.005 ;
        RECT 13.365 34.395 13.535 34.565 ;
        RECT 13.365 28.955 13.535 29.125 ;
        RECT 13.365 23.515 13.535 23.685 ;
        RECT 13.365 18.075 13.535 18.245 ;
        RECT 13.365 12.635 13.535 12.805 ;
        RECT 13.825 56.155 13.995 56.325 ;
        RECT 13.825 50.715 13.995 50.885 ;
        RECT 13.825 45.275 13.995 45.445 ;
        RECT 13.825 39.835 13.995 40.005 ;
        RECT 13.825 34.395 13.995 34.565 ;
        RECT 13.825 28.955 13.995 29.125 ;
        RECT 13.825 23.515 13.995 23.685 ;
        RECT 13.825 18.075 13.995 18.245 ;
        RECT 13.825 12.635 13.995 12.805 ;
        RECT 14.285 56.155 14.455 56.325 ;
        RECT 14.285 50.715 14.455 50.885 ;
        RECT 14.285 45.275 14.455 45.445 ;
        RECT 14.285 39.835 14.455 40.005 ;
        RECT 14.285 34.395 14.455 34.565 ;
        RECT 14.285 28.955 14.455 29.125 ;
        RECT 14.285 23.515 14.455 23.685 ;
        RECT 14.285 18.075 14.455 18.245 ;
        RECT 14.285 12.635 14.455 12.805 ;
        RECT 14.745 56.155 14.915 56.325 ;
        RECT 14.745 50.715 14.915 50.885 ;
        RECT 14.745 45.275 14.915 45.445 ;
        RECT 14.745 39.835 14.915 40.005 ;
        RECT 14.745 34.395 14.915 34.565 ;
        RECT 14.745 28.955 14.915 29.125 ;
        RECT 14.745 23.515 14.915 23.685 ;
        RECT 14.745 18.075 14.915 18.245 ;
        RECT 14.745 12.635 14.915 12.805 ;
        RECT 15.205 56.155 15.375 56.325 ;
        RECT 15.205 50.715 15.375 50.885 ;
        RECT 15.205 45.275 15.375 45.445 ;
        RECT 15.205 39.835 15.375 40.005 ;
        RECT 15.205 34.395 15.375 34.565 ;
        RECT 15.205 28.955 15.375 29.125 ;
        RECT 15.205 23.515 15.375 23.685 ;
        RECT 15.205 18.075 15.375 18.245 ;
        RECT 15.205 12.635 15.375 12.805 ;
        RECT 15.665 56.155 15.835 56.325 ;
        RECT 15.665 50.715 15.835 50.885 ;
        RECT 15.665 45.275 15.835 45.445 ;
        RECT 15.665 39.835 15.835 40.005 ;
        RECT 15.665 34.395 15.835 34.565 ;
        RECT 15.665 28.955 15.835 29.125 ;
        RECT 15.665 23.515 15.835 23.685 ;
        RECT 15.665 18.075 15.835 18.245 ;
        RECT 15.665 12.635 15.835 12.805 ;
        RECT 16.125 56.155 16.295 56.325 ;
        RECT 16.125 50.715 16.295 50.885 ;
        RECT 16.125 45.275 16.295 45.445 ;
        RECT 16.125 39.835 16.295 40.005 ;
        RECT 16.125 34.395 16.295 34.565 ;
        RECT 16.125 28.955 16.295 29.125 ;
        RECT 16.125 23.515 16.295 23.685 ;
        RECT 16.125 18.075 16.295 18.245 ;
        RECT 16.125 12.635 16.295 12.805 ;
        RECT 16.585 56.155 16.755 56.325 ;
        RECT 16.585 50.715 16.755 50.885 ;
        RECT 16.585 45.275 16.755 45.445 ;
        RECT 16.585 39.835 16.755 40.005 ;
        RECT 16.585 34.395 16.755 34.565 ;
        RECT 16.585 28.955 16.755 29.125 ;
        RECT 16.585 23.515 16.755 23.685 ;
        RECT 16.585 18.075 16.755 18.245 ;
        RECT 16.585 12.635 16.755 12.805 ;
        RECT 17.045 56.155 17.215 56.325 ;
        RECT 17.045 50.715 17.215 50.885 ;
        RECT 17.045 45.275 17.215 45.445 ;
        RECT 17.045 39.835 17.215 40.005 ;
        RECT 17.045 34.395 17.215 34.565 ;
        RECT 17.045 28.955 17.215 29.125 ;
        RECT 17.045 23.515 17.215 23.685 ;
        RECT 17.045 18.075 17.215 18.245 ;
        RECT 17.045 12.635 17.215 12.805 ;
        RECT 17.505 56.155 17.675 56.325 ;
        RECT 17.505 50.715 17.675 50.885 ;
        RECT 17.505 45.275 17.675 45.445 ;
        RECT 17.505 39.835 17.675 40.005 ;
        RECT 17.505 34.395 17.675 34.565 ;
        RECT 17.505 28.955 17.675 29.125 ;
        RECT 17.505 23.515 17.675 23.685 ;
        RECT 17.505 18.075 17.675 18.245 ;
        RECT 17.505 12.635 17.675 12.805 ;
        RECT 17.965 56.155 18.135 56.325 ;
        RECT 17.965 50.715 18.135 50.885 ;
        RECT 17.965 45.275 18.135 45.445 ;
        RECT 17.965 39.835 18.135 40.005 ;
        RECT 17.965 34.395 18.135 34.565 ;
        RECT 17.965 28.955 18.135 29.125 ;
        RECT 17.965 23.515 18.135 23.685 ;
        RECT 17.965 18.075 18.135 18.245 ;
        RECT 17.965 12.635 18.135 12.805 ;
        RECT 18.425 56.155 18.595 56.325 ;
        RECT 18.425 50.715 18.595 50.885 ;
        RECT 18.425 45.275 18.595 45.445 ;
        RECT 18.425 39.835 18.595 40.005 ;
        RECT 18.425 34.395 18.595 34.565 ;
        RECT 18.425 28.955 18.595 29.125 ;
        RECT 18.425 23.515 18.595 23.685 ;
        RECT 18.425 18.075 18.595 18.245 ;
        RECT 18.425 12.635 18.595 12.805 ;
        RECT 18.885 56.155 19.055 56.325 ;
        RECT 18.885 50.715 19.055 50.885 ;
        RECT 18.885 45.275 19.055 45.445 ;
        RECT 18.885 39.835 19.055 40.005 ;
        RECT 18.885 34.395 19.055 34.565 ;
        RECT 18.885 28.955 19.055 29.125 ;
        RECT 18.885 23.515 19.055 23.685 ;
        RECT 18.885 18.075 19.055 18.245 ;
        RECT 18.885 12.635 19.055 12.805 ;
        RECT 19.345 56.155 19.515 56.325 ;
        RECT 19.345 50.715 19.515 50.885 ;
        RECT 19.345 45.275 19.515 45.445 ;
        RECT 19.345 39.835 19.515 40.005 ;
        RECT 19.345 34.395 19.515 34.565 ;
        RECT 19.345 28.955 19.515 29.125 ;
        RECT 19.345 23.515 19.515 23.685 ;
        RECT 19.345 18.075 19.515 18.245 ;
        RECT 19.345 12.635 19.515 12.805 ;
        RECT 19.805 56.155 19.975 56.325 ;
        RECT 19.805 50.715 19.975 50.885 ;
        RECT 19.805 45.275 19.975 45.445 ;
        RECT 19.805 39.835 19.975 40.005 ;
        RECT 19.805 34.395 19.975 34.565 ;
        RECT 19.805 28.955 19.975 29.125 ;
        RECT 19.805 23.515 19.975 23.685 ;
        RECT 19.805 18.075 19.975 18.245 ;
        RECT 19.805 12.635 19.975 12.805 ;
        RECT 20.265 56.155 20.435 56.325 ;
        RECT 20.265 50.715 20.435 50.885 ;
        RECT 20.265 45.275 20.435 45.445 ;
        RECT 20.265 39.835 20.435 40.005 ;
        RECT 20.265 34.395 20.435 34.565 ;
        RECT 20.265 28.955 20.435 29.125 ;
        RECT 20.265 23.515 20.435 23.685 ;
        RECT 20.265 18.075 20.435 18.245 ;
        RECT 20.265 12.635 20.435 12.805 ;
        RECT 20.725 56.155 20.895 56.325 ;
        RECT 20.725 50.715 20.895 50.885 ;
        RECT 20.725 45.275 20.895 45.445 ;
        RECT 20.725 39.835 20.895 40.005 ;
        RECT 20.725 34.395 20.895 34.565 ;
        RECT 20.725 28.955 20.895 29.125 ;
        RECT 20.725 23.515 20.895 23.685 ;
        RECT 20.725 18.075 20.895 18.245 ;
        RECT 20.725 12.635 20.895 12.805 ;
        RECT 21.185 56.155 21.355 56.325 ;
        RECT 21.185 50.715 21.355 50.885 ;
        RECT 21.185 45.275 21.355 45.445 ;
        RECT 21.185 39.835 21.355 40.005 ;
        RECT 21.185 34.395 21.355 34.565 ;
        RECT 21.185 28.955 21.355 29.125 ;
        RECT 21.185 23.515 21.355 23.685 ;
        RECT 21.185 18.075 21.355 18.245 ;
        RECT 21.185 12.635 21.355 12.805 ;
        RECT 21.645 56.155 21.815 56.325 ;
        RECT 21.645 50.715 21.815 50.885 ;
        RECT 21.645 45.275 21.815 45.445 ;
        RECT 21.645 39.835 21.815 40.005 ;
        RECT 21.645 34.395 21.815 34.565 ;
        RECT 21.645 28.955 21.815 29.125 ;
        RECT 21.645 23.515 21.815 23.685 ;
        RECT 21.645 18.075 21.815 18.245 ;
        RECT 21.645 12.635 21.815 12.805 ;
        RECT 22.105 56.155 22.275 56.325 ;
        RECT 22.105 50.715 22.275 50.885 ;
        RECT 22.105 45.275 22.275 45.445 ;
        RECT 22.105 39.835 22.275 40.005 ;
        RECT 22.105 34.395 22.275 34.565 ;
        RECT 22.105 28.955 22.275 29.125 ;
        RECT 22.105 23.515 22.275 23.685 ;
        RECT 22.105 18.075 22.275 18.245 ;
        RECT 22.105 12.635 22.275 12.805 ;
        RECT 22.565 56.155 22.735 56.325 ;
        RECT 22.565 50.715 22.735 50.885 ;
        RECT 22.565 45.275 22.735 45.445 ;
        RECT 22.565 39.835 22.735 40.005 ;
        RECT 22.565 34.395 22.735 34.565 ;
        RECT 22.565 28.955 22.735 29.125 ;
        RECT 22.565 23.515 22.735 23.685 ;
        RECT 22.565 18.075 22.735 18.245 ;
        RECT 22.565 12.635 22.735 12.805 ;
        RECT 23.025 56.155 23.195 56.325 ;
        RECT 23.025 50.715 23.195 50.885 ;
        RECT 23.025 45.275 23.195 45.445 ;
        RECT 23.025 39.835 23.195 40.005 ;
        RECT 23.025 34.395 23.195 34.565 ;
        RECT 23.025 28.955 23.195 29.125 ;
        RECT 23.025 23.515 23.195 23.685 ;
        RECT 23.025 18.075 23.195 18.245 ;
        RECT 23.025 12.635 23.195 12.805 ;
        RECT 23.485 56.155 23.655 56.325 ;
        RECT 23.485 50.715 23.655 50.885 ;
        RECT 23.485 45.275 23.655 45.445 ;
        RECT 23.485 39.835 23.655 40.005 ;
        RECT 23.485 34.395 23.655 34.565 ;
        RECT 23.485 28.955 23.655 29.125 ;
        RECT 23.485 23.515 23.655 23.685 ;
        RECT 23.485 18.075 23.655 18.245 ;
        RECT 23.485 12.635 23.655 12.805 ;
        RECT 23.945 56.155 24.115 56.325 ;
        RECT 23.945 50.715 24.115 50.885 ;
        RECT 23.945 45.275 24.115 45.445 ;
        RECT 23.945 39.835 24.115 40.005 ;
        RECT 23.945 34.395 24.115 34.565 ;
        RECT 23.945 28.955 24.115 29.125 ;
        RECT 23.945 23.515 24.115 23.685 ;
        RECT 23.945 18.075 24.115 18.245 ;
        RECT 23.945 12.635 24.115 12.805 ;
        RECT 24.405 56.155 24.575 56.325 ;
        RECT 24.405 50.715 24.575 50.885 ;
        RECT 24.405 45.275 24.575 45.445 ;
        RECT 24.405 39.835 24.575 40.005 ;
        RECT 24.405 34.395 24.575 34.565 ;
        RECT 24.405 28.955 24.575 29.125 ;
        RECT 24.405 23.515 24.575 23.685 ;
        RECT 24.405 18.075 24.575 18.245 ;
        RECT 24.405 12.635 24.575 12.805 ;
        RECT 24.865 56.155 25.035 56.325 ;
        RECT 24.865 50.715 25.035 50.885 ;
        RECT 24.865 45.275 25.035 45.445 ;
        RECT 24.865 39.835 25.035 40.005 ;
        RECT 24.865 34.395 25.035 34.565 ;
        RECT 24.865 28.955 25.035 29.125 ;
        RECT 24.865 23.515 25.035 23.685 ;
        RECT 24.865 18.075 25.035 18.245 ;
        RECT 24.865 12.635 25.035 12.805 ;
        RECT 25.325 56.155 25.495 56.325 ;
        RECT 25.325 50.715 25.495 50.885 ;
        RECT 25.325 45.275 25.495 45.445 ;
        RECT 25.325 39.835 25.495 40.005 ;
        RECT 25.325 34.395 25.495 34.565 ;
        RECT 25.325 28.955 25.495 29.125 ;
        RECT 25.325 23.515 25.495 23.685 ;
        RECT 25.325 18.075 25.495 18.245 ;
        RECT 25.325 12.635 25.495 12.805 ;
        RECT 25.785 56.155 25.955 56.325 ;
        RECT 25.785 50.715 25.955 50.885 ;
        RECT 25.785 45.275 25.955 45.445 ;
        RECT 25.785 39.835 25.955 40.005 ;
        RECT 25.785 34.395 25.955 34.565 ;
        RECT 25.785 28.955 25.955 29.125 ;
        RECT 25.785 23.515 25.955 23.685 ;
        RECT 25.785 18.075 25.955 18.245 ;
        RECT 25.785 12.635 25.955 12.805 ;
        RECT 26.245 56.155 26.415 56.325 ;
        RECT 26.245 50.715 26.415 50.885 ;
        RECT 26.245 45.275 26.415 45.445 ;
        RECT 26.245 39.835 26.415 40.005 ;
        RECT 26.245 34.395 26.415 34.565 ;
        RECT 26.245 28.955 26.415 29.125 ;
        RECT 26.245 23.515 26.415 23.685 ;
        RECT 26.245 18.075 26.415 18.245 ;
        RECT 26.245 12.635 26.415 12.805 ;
        RECT 26.705 56.155 26.875 56.325 ;
        RECT 26.705 50.715 26.875 50.885 ;
        RECT 26.705 45.275 26.875 45.445 ;
        RECT 26.705 39.835 26.875 40.005 ;
        RECT 26.705 34.395 26.875 34.565 ;
        RECT 26.705 28.955 26.875 29.125 ;
        RECT 26.705 23.515 26.875 23.685 ;
        RECT 26.705 18.075 26.875 18.245 ;
        RECT 26.705 12.635 26.875 12.805 ;
        RECT 27.165 56.155 27.335 56.325 ;
        RECT 27.165 50.715 27.335 50.885 ;
        RECT 27.165 45.275 27.335 45.445 ;
        RECT 27.165 39.835 27.335 40.005 ;
        RECT 27.165 34.395 27.335 34.565 ;
        RECT 27.165 28.955 27.335 29.125 ;
        RECT 27.165 23.515 27.335 23.685 ;
        RECT 27.165 18.075 27.335 18.245 ;
        RECT 27.165 12.635 27.335 12.805 ;
        RECT 27.625 56.155 27.795 56.325 ;
        RECT 27.625 50.715 27.795 50.885 ;
        RECT 27.625 45.275 27.795 45.445 ;
        RECT 27.625 39.835 27.795 40.005 ;
        RECT 27.625 34.395 27.795 34.565 ;
        RECT 27.625 28.955 27.795 29.125 ;
        RECT 27.625 23.515 27.795 23.685 ;
        RECT 27.625 18.075 27.795 18.245 ;
        RECT 27.625 12.635 27.795 12.805 ;
        RECT 28.085 56.155 28.255 56.325 ;
        RECT 28.085 50.715 28.255 50.885 ;
        RECT 28.085 45.275 28.255 45.445 ;
        RECT 28.085 39.835 28.255 40.005 ;
        RECT 28.085 34.395 28.255 34.565 ;
        RECT 28.085 28.955 28.255 29.125 ;
        RECT 28.085 23.515 28.255 23.685 ;
        RECT 28.085 18.075 28.255 18.245 ;
        RECT 28.085 12.635 28.255 12.805 ;
        RECT 28.545 56.155 28.715 56.325 ;
        RECT 28.545 50.715 28.715 50.885 ;
        RECT 28.545 45.275 28.715 45.445 ;
        RECT 28.545 39.835 28.715 40.005 ;
        RECT 28.545 34.395 28.715 34.565 ;
        RECT 28.545 28.955 28.715 29.125 ;
        RECT 28.545 23.515 28.715 23.685 ;
        RECT 28.545 18.075 28.715 18.245 ;
        RECT 28.545 12.635 28.715 12.805 ;
        RECT 29.005 56.155 29.175 56.325 ;
        RECT 29.005 50.715 29.175 50.885 ;
        RECT 29.005 45.275 29.175 45.445 ;
        RECT 29.005 39.835 29.175 40.005 ;
        RECT 29.005 34.395 29.175 34.565 ;
        RECT 29.005 28.955 29.175 29.125 ;
        RECT 29.005 23.515 29.175 23.685 ;
        RECT 29.005 18.075 29.175 18.245 ;
        RECT 29.005 12.635 29.175 12.805 ;
        RECT 29.465 56.155 29.635 56.325 ;
        RECT 29.465 50.715 29.635 50.885 ;
        RECT 29.465 45.275 29.635 45.445 ;
        RECT 29.465 39.835 29.635 40.005 ;
        RECT 29.465 34.395 29.635 34.565 ;
        RECT 29.465 28.955 29.635 29.125 ;
        RECT 29.465 23.515 29.635 23.685 ;
        RECT 29.465 18.075 29.635 18.245 ;
        RECT 29.465 12.635 29.635 12.805 ;
        RECT 29.925 56.155 30.095 56.325 ;
        RECT 29.925 50.715 30.095 50.885 ;
        RECT 29.925 45.275 30.095 45.445 ;
        RECT 29.925 39.835 30.095 40.005 ;
        RECT 29.925 34.395 30.095 34.565 ;
        RECT 29.925 28.955 30.095 29.125 ;
        RECT 29.925 23.515 30.095 23.685 ;
        RECT 29.925 18.075 30.095 18.245 ;
        RECT 29.925 12.635 30.095 12.805 ;
        RECT 30.385 56.155 30.555 56.325 ;
        RECT 30.385 50.715 30.555 50.885 ;
        RECT 30.385 45.275 30.555 45.445 ;
        RECT 30.385 39.835 30.555 40.005 ;
        RECT 30.385 34.395 30.555 34.565 ;
        RECT 30.385 28.955 30.555 29.125 ;
        RECT 30.385 23.515 30.555 23.685 ;
        RECT 30.385 18.075 30.555 18.245 ;
        RECT 30.385 12.635 30.555 12.805 ;
        RECT 30.845 56.155 31.015 56.325 ;
        RECT 30.845 50.715 31.015 50.885 ;
        RECT 30.845 45.275 31.015 45.445 ;
        RECT 30.845 39.835 31.015 40.005 ;
        RECT 30.845 34.395 31.015 34.565 ;
        RECT 30.845 28.955 31.015 29.125 ;
        RECT 30.845 23.515 31.015 23.685 ;
        RECT 30.845 18.075 31.015 18.245 ;
        RECT 30.845 12.635 31.015 12.805 ;
        RECT 31.305 56.155 31.475 56.325 ;
        RECT 31.305 50.715 31.475 50.885 ;
        RECT 31.305 45.275 31.475 45.445 ;
        RECT 31.305 39.835 31.475 40.005 ;
        RECT 31.305 34.395 31.475 34.565 ;
        RECT 31.305 28.955 31.475 29.125 ;
        RECT 31.305 23.515 31.475 23.685 ;
        RECT 31.305 18.075 31.475 18.245 ;
        RECT 31.305 12.635 31.475 12.805 ;
        RECT 31.765 56.155 31.935 56.325 ;
        RECT 31.765 50.715 31.935 50.885 ;
        RECT 31.765 45.275 31.935 45.445 ;
        RECT 31.765 39.835 31.935 40.005 ;
        RECT 31.765 34.395 31.935 34.565 ;
        RECT 31.765 28.955 31.935 29.125 ;
        RECT 31.765 23.515 31.935 23.685 ;
        RECT 31.765 18.075 31.935 18.245 ;
        RECT 31.765 12.635 31.935 12.805 ;
        RECT 32.225 56.155 32.395 56.325 ;
        RECT 32.225 50.715 32.395 50.885 ;
        RECT 32.225 45.275 32.395 45.445 ;
        RECT 32.225 39.835 32.395 40.005 ;
        RECT 32.225 34.395 32.395 34.565 ;
        RECT 32.225 28.955 32.395 29.125 ;
        RECT 32.225 23.515 32.395 23.685 ;
        RECT 32.225 18.075 32.395 18.245 ;
        RECT 32.225 12.635 32.395 12.805 ;
        RECT 32.685 56.155 32.855 56.325 ;
        RECT 32.685 50.715 32.855 50.885 ;
        RECT 32.685 45.275 32.855 45.445 ;
        RECT 32.685 39.835 32.855 40.005 ;
        RECT 32.685 34.395 32.855 34.565 ;
        RECT 32.685 28.955 32.855 29.125 ;
        RECT 32.685 23.515 32.855 23.685 ;
        RECT 32.685 18.075 32.855 18.245 ;
        RECT 32.685 12.635 32.855 12.805 ;
        RECT 33.145 56.155 33.315 56.325 ;
        RECT 33.145 50.715 33.315 50.885 ;
        RECT 33.145 45.275 33.315 45.445 ;
        RECT 33.145 39.835 33.315 40.005 ;
        RECT 33.145 34.395 33.315 34.565 ;
        RECT 33.145 28.955 33.315 29.125 ;
        RECT 33.145 23.515 33.315 23.685 ;
        RECT 33.145 18.075 33.315 18.245 ;
        RECT 33.145 12.635 33.315 12.805 ;
        RECT 33.605 56.155 33.775 56.325 ;
        RECT 33.605 50.715 33.775 50.885 ;
        RECT 33.605 45.275 33.775 45.445 ;
        RECT 33.605 39.835 33.775 40.005 ;
        RECT 33.605 34.395 33.775 34.565 ;
        RECT 33.605 28.955 33.775 29.125 ;
        RECT 33.605 23.515 33.775 23.685 ;
        RECT 33.605 18.075 33.775 18.245 ;
        RECT 33.605 12.635 33.775 12.805 ;
        RECT 34.065 56.155 34.235 56.325 ;
        RECT 34.065 50.715 34.235 50.885 ;
        RECT 34.065 45.275 34.235 45.445 ;
        RECT 34.065 39.835 34.235 40.005 ;
        RECT 34.065 34.395 34.235 34.565 ;
        RECT 34.065 28.955 34.235 29.125 ;
        RECT 34.065 23.515 34.235 23.685 ;
        RECT 34.065 18.075 34.235 18.245 ;
        RECT 34.065 12.635 34.235 12.805 ;
        RECT 34.525 56.155 34.695 56.325 ;
        RECT 34.525 50.715 34.695 50.885 ;
        RECT 34.525 45.275 34.695 45.445 ;
        RECT 34.525 39.835 34.695 40.005 ;
        RECT 34.525 34.395 34.695 34.565 ;
        RECT 34.525 28.955 34.695 29.125 ;
        RECT 34.525 23.515 34.695 23.685 ;
        RECT 34.525 18.075 34.695 18.245 ;
        RECT 34.525 12.635 34.695 12.805 ;
        RECT 34.985 56.155 35.155 56.325 ;
        RECT 34.985 50.715 35.155 50.885 ;
        RECT 34.985 45.275 35.155 45.445 ;
        RECT 34.985 39.835 35.155 40.005 ;
        RECT 34.985 34.395 35.155 34.565 ;
        RECT 34.985 28.955 35.155 29.125 ;
        RECT 34.985 23.515 35.155 23.685 ;
        RECT 34.985 18.075 35.155 18.245 ;
        RECT 34.985 12.635 35.155 12.805 ;
        RECT 35.445 56.155 35.615 56.325 ;
        RECT 35.445 50.715 35.615 50.885 ;
        RECT 35.445 45.275 35.615 45.445 ;
        RECT 35.445 39.835 35.615 40.005 ;
        RECT 35.445 34.395 35.615 34.565 ;
        RECT 35.445 28.955 35.615 29.125 ;
        RECT 35.445 23.515 35.615 23.685 ;
        RECT 35.445 18.075 35.615 18.245 ;
        RECT 35.445 12.635 35.615 12.805 ;
        RECT 35.905 56.155 36.075 56.325 ;
        RECT 35.905 50.715 36.075 50.885 ;
        RECT 35.905 45.275 36.075 45.445 ;
        RECT 35.905 39.835 36.075 40.005 ;
        RECT 35.905 34.395 36.075 34.565 ;
        RECT 35.905 28.955 36.075 29.125 ;
        RECT 35.905 23.515 36.075 23.685 ;
        RECT 35.905 18.075 36.075 18.245 ;
        RECT 35.905 12.635 36.075 12.805 ;
        RECT 36.365 56.155 36.535 56.325 ;
        RECT 36.365 50.715 36.535 50.885 ;
        RECT 36.365 45.275 36.535 45.445 ;
        RECT 36.365 39.835 36.535 40.005 ;
        RECT 36.365 34.395 36.535 34.565 ;
        RECT 36.365 28.955 36.535 29.125 ;
        RECT 36.365 23.515 36.535 23.685 ;
        RECT 36.365 18.075 36.535 18.245 ;
        RECT 36.365 12.635 36.535 12.805 ;
        RECT 36.825 56.155 36.995 56.325 ;
        RECT 36.825 50.715 36.995 50.885 ;
        RECT 36.825 45.275 36.995 45.445 ;
        RECT 36.825 39.835 36.995 40.005 ;
        RECT 36.825 34.395 36.995 34.565 ;
        RECT 36.825 28.955 36.995 29.125 ;
        RECT 36.825 23.515 36.995 23.685 ;
        RECT 36.825 18.075 36.995 18.245 ;
        RECT 36.825 12.635 36.995 12.805 ;
        RECT 37.285 56.155 37.455 56.325 ;
        RECT 37.285 50.715 37.455 50.885 ;
        RECT 37.285 45.275 37.455 45.445 ;
        RECT 37.285 39.835 37.455 40.005 ;
        RECT 37.285 34.395 37.455 34.565 ;
        RECT 37.285 28.955 37.455 29.125 ;
        RECT 37.285 23.515 37.455 23.685 ;
        RECT 37.285 18.075 37.455 18.245 ;
        RECT 37.285 12.635 37.455 12.805 ;
        RECT 37.745 56.155 37.915 56.325 ;
        RECT 37.745 50.715 37.915 50.885 ;
        RECT 37.745 45.275 37.915 45.445 ;
        RECT 37.745 39.835 37.915 40.005 ;
        RECT 37.745 34.395 37.915 34.565 ;
        RECT 37.745 28.955 37.915 29.125 ;
        RECT 37.745 23.515 37.915 23.685 ;
        RECT 37.745 18.075 37.915 18.245 ;
        RECT 37.745 12.635 37.915 12.805 ;
        RECT 38.205 56.155 38.375 56.325 ;
        RECT 38.205 50.715 38.375 50.885 ;
        RECT 38.205 45.275 38.375 45.445 ;
        RECT 38.205 39.835 38.375 40.005 ;
        RECT 38.205 34.395 38.375 34.565 ;
        RECT 38.205 28.955 38.375 29.125 ;
        RECT 38.205 23.515 38.375 23.685 ;
        RECT 38.205 18.075 38.375 18.245 ;
        RECT 38.205 12.635 38.375 12.805 ;
        RECT 38.665 56.155 38.835 56.325 ;
        RECT 38.665 50.715 38.835 50.885 ;
        RECT 38.665 45.275 38.835 45.445 ;
        RECT 38.665 39.835 38.835 40.005 ;
        RECT 38.665 34.395 38.835 34.565 ;
        RECT 38.665 28.955 38.835 29.125 ;
        RECT 38.665 23.515 38.835 23.685 ;
        RECT 38.665 18.075 38.835 18.245 ;
        RECT 38.665 12.635 38.835 12.805 ;
        RECT 39.125 56.155 39.295 56.325 ;
        RECT 39.125 50.715 39.295 50.885 ;
        RECT 39.125 45.275 39.295 45.445 ;
        RECT 39.125 39.835 39.295 40.005 ;
        RECT 39.125 34.395 39.295 34.565 ;
        RECT 39.125 28.955 39.295 29.125 ;
        RECT 39.125 23.515 39.295 23.685 ;
        RECT 39.125 18.075 39.295 18.245 ;
        RECT 39.125 12.635 39.295 12.805 ;
        RECT 39.585 56.155 39.755 56.325 ;
        RECT 39.585 50.715 39.755 50.885 ;
        RECT 39.585 45.275 39.755 45.445 ;
        RECT 39.585 39.835 39.755 40.005 ;
        RECT 39.585 34.395 39.755 34.565 ;
        RECT 39.585 28.955 39.755 29.125 ;
        RECT 39.585 23.515 39.755 23.685 ;
        RECT 39.585 18.075 39.755 18.245 ;
        RECT 39.585 12.635 39.755 12.805 ;
        RECT 40.045 56.155 40.215 56.325 ;
        RECT 40.045 50.715 40.215 50.885 ;
        RECT 40.045 45.275 40.215 45.445 ;
        RECT 40.045 39.835 40.215 40.005 ;
        RECT 40.045 34.395 40.215 34.565 ;
        RECT 40.045 28.955 40.215 29.125 ;
        RECT 40.045 23.515 40.215 23.685 ;
        RECT 40.045 18.075 40.215 18.245 ;
        RECT 40.045 12.635 40.215 12.805 ;
        RECT 40.505 56.155 40.675 56.325 ;
        RECT 40.505 50.715 40.675 50.885 ;
        RECT 40.505 45.275 40.675 45.445 ;
        RECT 40.505 39.835 40.675 40.005 ;
        RECT 40.505 34.395 40.675 34.565 ;
        RECT 40.505 28.955 40.675 29.125 ;
        RECT 40.505 23.515 40.675 23.685 ;
        RECT 40.505 18.075 40.675 18.245 ;
        RECT 40.505 12.635 40.675 12.805 ;
        RECT 40.965 56.155 41.135 56.325 ;
        RECT 40.965 50.715 41.135 50.885 ;
        RECT 40.965 45.275 41.135 45.445 ;
        RECT 40.965 39.835 41.135 40.005 ;
        RECT 40.965 34.395 41.135 34.565 ;
        RECT 40.965 28.955 41.135 29.125 ;
        RECT 40.965 23.515 41.135 23.685 ;
        RECT 40.965 18.075 41.135 18.245 ;
        RECT 40.965 12.635 41.135 12.805 ;
        RECT 41.425 56.155 41.595 56.325 ;
        RECT 41.425 50.715 41.595 50.885 ;
        RECT 41.425 45.275 41.595 45.445 ;
        RECT 41.425 39.835 41.595 40.005 ;
        RECT 41.425 34.395 41.595 34.565 ;
        RECT 41.425 28.955 41.595 29.125 ;
        RECT 41.425 23.515 41.595 23.685 ;
        RECT 41.425 18.075 41.595 18.245 ;
        RECT 41.425 12.635 41.595 12.805 ;
        RECT 41.885 56.155 42.055 56.325 ;
        RECT 41.885 50.715 42.055 50.885 ;
        RECT 41.885 45.275 42.055 45.445 ;
        RECT 41.885 39.835 42.055 40.005 ;
        RECT 41.885 34.395 42.055 34.565 ;
        RECT 41.885 28.955 42.055 29.125 ;
        RECT 41.885 23.515 42.055 23.685 ;
        RECT 41.885 18.075 42.055 18.245 ;
        RECT 41.885 12.635 42.055 12.805 ;
        RECT 42.345 56.155 42.515 56.325 ;
        RECT 42.345 50.715 42.515 50.885 ;
        RECT 42.345 45.275 42.515 45.445 ;
        RECT 42.345 39.835 42.515 40.005 ;
        RECT 42.345 34.395 42.515 34.565 ;
        RECT 42.345 28.955 42.515 29.125 ;
        RECT 42.345 23.515 42.515 23.685 ;
        RECT 42.345 18.075 42.515 18.245 ;
        RECT 42.345 12.635 42.515 12.805 ;
        RECT 42.805 56.155 42.975 56.325 ;
        RECT 42.805 50.715 42.975 50.885 ;
        RECT 42.805 45.275 42.975 45.445 ;
        RECT 42.805 39.835 42.975 40.005 ;
        RECT 42.805 34.395 42.975 34.565 ;
        RECT 42.805 28.955 42.975 29.125 ;
        RECT 42.805 23.515 42.975 23.685 ;
        RECT 42.805 18.075 42.975 18.245 ;
        RECT 42.805 12.635 42.975 12.805 ;
        RECT 43.265 56.155 43.435 56.325 ;
        RECT 43.265 50.715 43.435 50.885 ;
        RECT 43.265 45.275 43.435 45.445 ;
        RECT 43.265 39.835 43.435 40.005 ;
        RECT 43.265 34.395 43.435 34.565 ;
        RECT 43.265 28.955 43.435 29.125 ;
        RECT 43.265 23.515 43.435 23.685 ;
        RECT 43.265 18.075 43.435 18.245 ;
        RECT 43.265 12.635 43.435 12.805 ;
        RECT 43.725 56.155 43.895 56.325 ;
        RECT 43.725 50.715 43.895 50.885 ;
        RECT 43.725 45.275 43.895 45.445 ;
        RECT 43.725 39.835 43.895 40.005 ;
        RECT 43.725 34.395 43.895 34.565 ;
        RECT 43.725 28.955 43.895 29.125 ;
        RECT 43.725 23.515 43.895 23.685 ;
        RECT 43.725 18.075 43.895 18.245 ;
        RECT 43.725 12.635 43.895 12.805 ;
        RECT 44.185 56.155 44.355 56.325 ;
        RECT 44.185 50.715 44.355 50.885 ;
        RECT 44.185 45.275 44.355 45.445 ;
        RECT 44.185 39.835 44.355 40.005 ;
        RECT 44.185 34.395 44.355 34.565 ;
        RECT 44.185 28.955 44.355 29.125 ;
        RECT 44.185 23.515 44.355 23.685 ;
        RECT 44.185 18.075 44.355 18.245 ;
        RECT 44.185 12.635 44.355 12.805 ;
        RECT 44.645 56.155 44.815 56.325 ;
        RECT 44.645 50.715 44.815 50.885 ;
        RECT 44.645 45.275 44.815 45.445 ;
        RECT 44.645 39.835 44.815 40.005 ;
        RECT 44.645 34.395 44.815 34.565 ;
        RECT 44.645 28.955 44.815 29.125 ;
        RECT 44.645 23.515 44.815 23.685 ;
        RECT 44.645 18.075 44.815 18.245 ;
        RECT 44.645 12.635 44.815 12.805 ;
        RECT 45.105 56.155 45.275 56.325 ;
        RECT 45.105 50.715 45.275 50.885 ;
        RECT 45.105 45.275 45.275 45.445 ;
        RECT 45.105 39.835 45.275 40.005 ;
        RECT 45.105 34.395 45.275 34.565 ;
        RECT 45.105 28.955 45.275 29.125 ;
        RECT 45.105 23.515 45.275 23.685 ;
        RECT 45.105 18.075 45.275 18.245 ;
        RECT 45.105 12.635 45.275 12.805 ;
        RECT 45.565 56.155 45.735 56.325 ;
        RECT 45.565 50.715 45.735 50.885 ;
        RECT 45.565 45.275 45.735 45.445 ;
        RECT 45.565 39.835 45.735 40.005 ;
        RECT 45.565 34.395 45.735 34.565 ;
        RECT 45.565 28.955 45.735 29.125 ;
        RECT 45.565 23.515 45.735 23.685 ;
        RECT 45.565 18.075 45.735 18.245 ;
        RECT 45.565 12.635 45.735 12.805 ;
        RECT 46.025 56.155 46.195 56.325 ;
        RECT 46.025 50.715 46.195 50.885 ;
        RECT 46.025 45.275 46.195 45.445 ;
        RECT 46.025 39.835 46.195 40.005 ;
        RECT 46.025 34.395 46.195 34.565 ;
        RECT 46.025 28.955 46.195 29.125 ;
        RECT 46.025 23.515 46.195 23.685 ;
        RECT 46.025 18.075 46.195 18.245 ;
        RECT 46.025 12.635 46.195 12.805 ;
        RECT 46.485 56.155 46.655 56.325 ;
        RECT 46.485 50.715 46.655 50.885 ;
        RECT 46.485 45.275 46.655 45.445 ;
        RECT 46.485 39.835 46.655 40.005 ;
        RECT 46.485 34.395 46.655 34.565 ;
        RECT 46.485 28.955 46.655 29.125 ;
        RECT 46.485 23.515 46.655 23.685 ;
        RECT 46.485 18.075 46.655 18.245 ;
        RECT 46.485 12.635 46.655 12.805 ;
        RECT 46.945 56.155 47.115 56.325 ;
        RECT 46.945 50.715 47.115 50.885 ;
        RECT 46.945 45.275 47.115 45.445 ;
        RECT 46.945 39.835 47.115 40.005 ;
        RECT 46.945 34.395 47.115 34.565 ;
        RECT 46.945 28.955 47.115 29.125 ;
        RECT 46.945 23.515 47.115 23.685 ;
        RECT 46.945 18.075 47.115 18.245 ;
        RECT 46.945 12.635 47.115 12.805 ;
        RECT 47.405 56.155 47.575 56.325 ;
        RECT 47.405 50.715 47.575 50.885 ;
        RECT 47.405 45.275 47.575 45.445 ;
        RECT 47.405 39.835 47.575 40.005 ;
        RECT 47.405 34.395 47.575 34.565 ;
        RECT 47.405 28.955 47.575 29.125 ;
        RECT 47.405 23.515 47.575 23.685 ;
        RECT 47.405 18.075 47.575 18.245 ;
        RECT 47.405 12.635 47.575 12.805 ;
        RECT 47.865 56.155 48.035 56.325 ;
        RECT 47.865 50.715 48.035 50.885 ;
        RECT 47.865 45.275 48.035 45.445 ;
        RECT 47.865 39.835 48.035 40.005 ;
        RECT 47.865 34.395 48.035 34.565 ;
        RECT 47.865 28.955 48.035 29.125 ;
        RECT 47.865 23.515 48.035 23.685 ;
        RECT 47.865 18.075 48.035 18.245 ;
        RECT 47.865 12.635 48.035 12.805 ;
        RECT 48.325 56.155 48.495 56.325 ;
        RECT 48.325 50.715 48.495 50.885 ;
        RECT 48.325 45.275 48.495 45.445 ;
        RECT 48.325 39.835 48.495 40.005 ;
        RECT 48.325 34.395 48.495 34.565 ;
        RECT 48.325 28.955 48.495 29.125 ;
        RECT 48.325 23.515 48.495 23.685 ;
        RECT 48.325 18.075 48.495 18.245 ;
        RECT 48.325 12.635 48.495 12.805 ;
        RECT 48.785 56.155 48.955 56.325 ;
        RECT 48.785 50.715 48.955 50.885 ;
        RECT 48.785 45.275 48.955 45.445 ;
        RECT 48.785 39.835 48.955 40.005 ;
        RECT 48.785 34.395 48.955 34.565 ;
        RECT 48.785 28.955 48.955 29.125 ;
        RECT 48.785 23.515 48.955 23.685 ;
        RECT 48.785 18.075 48.955 18.245 ;
        RECT 48.785 12.635 48.955 12.805 ;
        RECT 49.245 56.155 49.415 56.325 ;
        RECT 49.245 50.715 49.415 50.885 ;
        RECT 49.245 45.275 49.415 45.445 ;
        RECT 49.245 39.835 49.415 40.005 ;
        RECT 49.245 34.395 49.415 34.565 ;
        RECT 49.245 28.955 49.415 29.125 ;
        RECT 49.245 23.515 49.415 23.685 ;
        RECT 49.245 18.075 49.415 18.245 ;
        RECT 49.245 12.635 49.415 12.805 ;
        RECT 49.705 56.155 49.875 56.325 ;
        RECT 49.705 50.715 49.875 50.885 ;
        RECT 49.705 45.275 49.875 45.445 ;
        RECT 49.705 39.835 49.875 40.005 ;
        RECT 49.705 34.395 49.875 34.565 ;
        RECT 49.705 28.955 49.875 29.125 ;
        RECT 49.705 23.515 49.875 23.685 ;
        RECT 49.705 18.075 49.875 18.245 ;
        RECT 49.705 12.635 49.875 12.805 ;
        RECT 50.165 56.155 50.335 56.325 ;
        RECT 50.165 50.715 50.335 50.885 ;
        RECT 50.165 45.275 50.335 45.445 ;
        RECT 50.165 39.835 50.335 40.005 ;
        RECT 50.165 34.395 50.335 34.565 ;
        RECT 50.165 28.955 50.335 29.125 ;
        RECT 50.165 23.515 50.335 23.685 ;
        RECT 50.165 18.075 50.335 18.245 ;
        RECT 50.165 12.635 50.335 12.805 ;
        RECT 50.625 56.155 50.795 56.325 ;
        RECT 50.625 50.715 50.795 50.885 ;
        RECT 50.625 45.275 50.795 45.445 ;
        RECT 50.625 39.835 50.795 40.005 ;
        RECT 50.625 34.395 50.795 34.565 ;
        RECT 50.625 28.955 50.795 29.125 ;
        RECT 50.625 23.515 50.795 23.685 ;
        RECT 50.625 18.075 50.795 18.245 ;
        RECT 50.625 12.635 50.795 12.805 ;
        RECT 51.085 56.155 51.255 56.325 ;
        RECT 51.085 50.715 51.255 50.885 ;
        RECT 51.085 45.275 51.255 45.445 ;
        RECT 51.085 39.835 51.255 40.005 ;
        RECT 51.085 34.395 51.255 34.565 ;
        RECT 51.085 28.955 51.255 29.125 ;
        RECT 51.085 23.515 51.255 23.685 ;
        RECT 51.085 18.075 51.255 18.245 ;
        RECT 51.085 12.635 51.255 12.805 ;
        RECT 51.545 56.155 51.715 56.325 ;
        RECT 51.545 50.715 51.715 50.885 ;
        RECT 51.545 45.275 51.715 45.445 ;
        RECT 51.545 39.835 51.715 40.005 ;
        RECT 51.545 34.395 51.715 34.565 ;
        RECT 51.545 28.955 51.715 29.125 ;
        RECT 51.545 23.515 51.715 23.685 ;
        RECT 51.545 18.075 51.715 18.245 ;
        RECT 51.545 12.635 51.715 12.805 ;
        RECT 52.005 56.155 52.175 56.325 ;
        RECT 52.005 50.715 52.175 50.885 ;
        RECT 52.005 45.275 52.175 45.445 ;
        RECT 52.005 39.835 52.175 40.005 ;
        RECT 52.005 34.395 52.175 34.565 ;
        RECT 52.005 28.955 52.175 29.125 ;
        RECT 52.005 23.515 52.175 23.685 ;
        RECT 52.005 18.075 52.175 18.245 ;
        RECT 52.005 12.635 52.175 12.805 ;
        RECT 52.465 56.155 52.635 56.325 ;
        RECT 52.465 50.715 52.635 50.885 ;
        RECT 52.465 45.275 52.635 45.445 ;
        RECT 52.465 39.835 52.635 40.005 ;
        RECT 52.465 34.395 52.635 34.565 ;
        RECT 52.465 28.955 52.635 29.125 ;
        RECT 52.465 23.515 52.635 23.685 ;
        RECT 52.465 18.075 52.635 18.245 ;
        RECT 52.465 12.635 52.635 12.805 ;
        RECT 52.925 56.155 53.095 56.325 ;
        RECT 52.925 50.715 53.095 50.885 ;
        RECT 52.925 45.275 53.095 45.445 ;
        RECT 52.925 39.835 53.095 40.005 ;
        RECT 52.925 34.395 53.095 34.565 ;
        RECT 52.925 28.955 53.095 29.125 ;
        RECT 52.925 23.515 53.095 23.685 ;
        RECT 52.925 18.075 53.095 18.245 ;
        RECT 52.925 12.635 53.095 12.805 ;
        RECT 53.385 56.155 53.555 56.325 ;
        RECT 53.385 50.715 53.555 50.885 ;
        RECT 53.385 45.275 53.555 45.445 ;
        RECT 53.385 39.835 53.555 40.005 ;
        RECT 53.385 34.395 53.555 34.565 ;
        RECT 53.385 28.955 53.555 29.125 ;
        RECT 53.385 23.515 53.555 23.685 ;
        RECT 53.385 18.075 53.555 18.245 ;
        RECT 53.385 12.635 53.555 12.805 ;
        RECT 53.845 56.155 54.015 56.325 ;
        RECT 53.845 50.715 54.015 50.885 ;
        RECT 53.845 45.275 54.015 45.445 ;
        RECT 53.845 39.835 54.015 40.005 ;
        RECT 53.845 34.395 54.015 34.565 ;
        RECT 53.845 28.955 54.015 29.125 ;
        RECT 53.845 23.515 54.015 23.685 ;
        RECT 53.845 18.075 54.015 18.245 ;
        RECT 53.845 12.635 54.015 12.805 ;
        RECT 54.305 56.155 54.475 56.325 ;
        RECT 54.305 50.715 54.475 50.885 ;
        RECT 54.305 45.275 54.475 45.445 ;
        RECT 54.305 39.835 54.475 40.005 ;
        RECT 54.305 34.395 54.475 34.565 ;
        RECT 54.305 28.955 54.475 29.125 ;
        RECT 54.305 23.515 54.475 23.685 ;
        RECT 54.305 18.075 54.475 18.245 ;
        RECT 54.305 12.635 54.475 12.805 ;
        RECT 54.765 56.155 54.935 56.325 ;
        RECT 54.765 50.715 54.935 50.885 ;
        RECT 54.765 45.275 54.935 45.445 ;
        RECT 54.765 39.835 54.935 40.005 ;
        RECT 54.765 34.395 54.935 34.565 ;
        RECT 54.765 28.955 54.935 29.125 ;
        RECT 54.765 23.515 54.935 23.685 ;
        RECT 54.765 18.075 54.935 18.245 ;
        RECT 54.765 12.635 54.935 12.805 ;
        RECT 55.225 56.155 55.395 56.325 ;
        RECT 55.225 50.715 55.395 50.885 ;
        RECT 55.225 45.275 55.395 45.445 ;
        RECT 55.225 39.835 55.395 40.005 ;
        RECT 55.225 34.395 55.395 34.565 ;
        RECT 55.225 28.955 55.395 29.125 ;
        RECT 55.225 23.515 55.395 23.685 ;
        RECT 55.225 18.075 55.395 18.245 ;
        RECT 55.225 12.635 55.395 12.805 ;
        RECT 55.685 56.155 55.855 56.325 ;
        RECT 55.685 50.715 55.855 50.885 ;
        RECT 55.685 45.275 55.855 45.445 ;
        RECT 55.685 39.835 55.855 40.005 ;
        RECT 55.685 34.395 55.855 34.565 ;
        RECT 55.685 28.955 55.855 29.125 ;
        RECT 55.685 23.515 55.855 23.685 ;
        RECT 55.685 18.075 55.855 18.245 ;
        RECT 55.685 12.635 55.855 12.805 ;
        RECT 56.145 56.155 56.315 56.325 ;
        RECT 56.145 50.715 56.315 50.885 ;
        RECT 56.145 45.275 56.315 45.445 ;
        RECT 56.145 39.835 56.315 40.005 ;
        RECT 56.145 34.395 56.315 34.565 ;
        RECT 56.145 28.955 56.315 29.125 ;
        RECT 56.145 23.515 56.315 23.685 ;
        RECT 56.145 18.075 56.315 18.245 ;
        RECT 56.145 12.635 56.315 12.805 ;
        RECT 56.605 56.155 56.775 56.325 ;
        RECT 56.605 50.715 56.775 50.885 ;
        RECT 56.605 45.275 56.775 45.445 ;
        RECT 56.605 39.835 56.775 40.005 ;
        RECT 56.605 34.395 56.775 34.565 ;
        RECT 56.605 28.955 56.775 29.125 ;
        RECT 56.605 23.515 56.775 23.685 ;
        RECT 56.605 18.075 56.775 18.245 ;
        RECT 56.605 12.635 56.775 12.805 ;
        RECT 57.065 56.155 57.235 56.325 ;
        RECT 57.065 50.715 57.235 50.885 ;
        RECT 57.065 45.275 57.235 45.445 ;
        RECT 57.065 39.835 57.235 40.005 ;
        RECT 57.065 34.395 57.235 34.565 ;
        RECT 57.065 28.955 57.235 29.125 ;
        RECT 57.065 23.515 57.235 23.685 ;
        RECT 57.065 18.075 57.235 18.245 ;
        RECT 57.065 12.635 57.235 12.805 ;
        RECT 57.525 56.155 57.695 56.325 ;
        RECT 57.525 50.715 57.695 50.885 ;
        RECT 57.525 45.275 57.695 45.445 ;
        RECT 57.525 39.835 57.695 40.005 ;
        RECT 57.525 34.395 57.695 34.565 ;
        RECT 57.525 28.955 57.695 29.125 ;
        RECT 57.525 23.515 57.695 23.685 ;
        RECT 57.525 18.075 57.695 18.245 ;
        RECT 57.525 12.635 57.695 12.805 ;
        RECT 57.985 56.155 58.155 56.325 ;
        RECT 57.985 50.715 58.155 50.885 ;
        RECT 57.985 45.275 58.155 45.445 ;
        RECT 57.985 39.835 58.155 40.005 ;
        RECT 57.985 34.395 58.155 34.565 ;
        RECT 57.985 28.955 58.155 29.125 ;
        RECT 57.985 23.515 58.155 23.685 ;
        RECT 57.985 18.075 58.155 18.245 ;
        RECT 57.985 12.635 58.155 12.805 ;
        RECT 58.445 56.155 58.615 56.325 ;
        RECT 58.445 50.715 58.615 50.885 ;
        RECT 58.445 45.275 58.615 45.445 ;
        RECT 58.445 39.835 58.615 40.005 ;
        RECT 58.445 34.395 58.615 34.565 ;
        RECT 58.445 28.955 58.615 29.125 ;
        RECT 58.445 23.515 58.615 23.685 ;
        RECT 58.445 18.075 58.615 18.245 ;
        RECT 58.445 12.635 58.615 12.805 ;
        RECT 58.905 56.155 59.075 56.325 ;
        RECT 58.905 50.715 59.075 50.885 ;
        RECT 58.905 45.275 59.075 45.445 ;
        RECT 58.905 39.835 59.075 40.005 ;
        RECT 58.905 34.395 59.075 34.565 ;
        RECT 58.905 28.955 59.075 29.125 ;
        RECT 58.905 23.515 59.075 23.685 ;
        RECT 58.905 18.075 59.075 18.245 ;
        RECT 58.905 12.635 59.075 12.805 ;
        RECT 59.365 56.155 59.535 56.325 ;
        RECT 59.365 50.715 59.535 50.885 ;
        RECT 59.365 45.275 59.535 45.445 ;
        RECT 59.365 39.835 59.535 40.005 ;
        RECT 59.365 34.395 59.535 34.565 ;
        RECT 59.365 28.955 59.535 29.125 ;
        RECT 59.365 23.515 59.535 23.685 ;
        RECT 59.365 18.075 59.535 18.245 ;
        RECT 59.365 12.635 59.535 12.805 ;
        RECT 59.825 56.155 59.995 56.325 ;
        RECT 59.825 50.715 59.995 50.885 ;
        RECT 59.825 45.275 59.995 45.445 ;
        RECT 59.825 39.835 59.995 40.005 ;
        RECT 59.825 34.395 59.995 34.565 ;
        RECT 59.825 28.955 59.995 29.125 ;
        RECT 59.825 23.515 59.995 23.685 ;
        RECT 59.825 18.075 59.995 18.245 ;
        RECT 59.825 12.635 59.995 12.805 ;
        RECT 60.285 56.155 60.455 56.325 ;
        RECT 60.285 50.715 60.455 50.885 ;
        RECT 60.285 45.275 60.455 45.445 ;
        RECT 60.285 39.835 60.455 40.005 ;
        RECT 60.285 34.395 60.455 34.565 ;
        RECT 60.285 28.955 60.455 29.125 ;
        RECT 60.285 23.515 60.455 23.685 ;
        RECT 60.285 18.075 60.455 18.245 ;
        RECT 60.285 12.635 60.455 12.805 ;
        RECT 60.745 56.155 60.915 56.325 ;
        RECT 60.745 50.715 60.915 50.885 ;
        RECT 60.745 45.275 60.915 45.445 ;
        RECT 60.745 39.835 60.915 40.005 ;
        RECT 60.745 34.395 60.915 34.565 ;
        RECT 60.745 28.955 60.915 29.125 ;
        RECT 60.745 23.515 60.915 23.685 ;
        RECT 60.745 18.075 60.915 18.245 ;
        RECT 60.745 12.635 60.915 12.805 ;
        RECT 61.205 56.155 61.375 56.325 ;
      LAYER via2 ;
        RECT 11.05 56.48 11.25 56.68 ;
        RECT 11.05 52.4 11.25 52.6 ;
        RECT 11.05 48.32 11.25 48.52 ;
        RECT 11.05 44.24 11.25 44.44 ;
        RECT 11.05 40.16 11.25 40.36 ;
        RECT 11.05 36.08 11.25 36.28 ;
        RECT 11.05 32 11.25 32.2 ;
        RECT 11.05 27.92 11.25 28.12 ;
        RECT 11.05 23.84 11.25 24.04 ;
        RECT 11.05 19.76 11.25 19.96 ;
        RECT 11.05 15.68 11.25 15.88 ;
        RECT 11.05 11.6 11.25 11.8 ;
        RECT 13.81 56.48 14.01 56.68 ;
        RECT 13.81 52.4 14.01 52.6 ;
        RECT 13.81 48.32 14.01 48.52 ;
        RECT 13.81 44.24 14.01 44.44 ;
        RECT 13.81 40.16 14.01 40.36 ;
        RECT 13.81 36.08 14.01 36.28 ;
        RECT 13.81 32 14.01 32.2 ;
        RECT 13.81 27.92 14.01 28.12 ;
        RECT 13.81 23.84 14.01 24.04 ;
        RECT 13.81 19.76 14.01 19.96 ;
        RECT 13.81 15.68 14.01 15.88 ;
        RECT 13.81 11.6 14.01 11.8 ;
        RECT 16.57 56.48 16.77 56.68 ;
        RECT 16.57 52.4 16.77 52.6 ;
        RECT 16.57 48.32 16.77 48.52 ;
        RECT 16.57 44.24 16.77 44.44 ;
        RECT 16.57 40.16 16.77 40.36 ;
        RECT 16.57 36.08 16.77 36.28 ;
        RECT 16.57 32 16.77 32.2 ;
        RECT 16.57 27.92 16.77 28.12 ;
        RECT 16.57 23.84 16.77 24.04 ;
        RECT 16.57 19.76 16.77 19.96 ;
        RECT 16.57 15.68 16.77 15.88 ;
        RECT 16.57 11.6 16.77 11.8 ;
        RECT 19.33 56.48 19.53 56.68 ;
        RECT 19.33 52.4 19.53 52.6 ;
        RECT 19.33 48.32 19.53 48.52 ;
        RECT 19.33 44.24 19.53 44.44 ;
        RECT 19.33 40.16 19.53 40.36 ;
        RECT 19.33 36.08 19.53 36.28 ;
        RECT 19.33 32 19.53 32.2 ;
        RECT 19.33 27.92 19.53 28.12 ;
        RECT 19.33 23.84 19.53 24.04 ;
        RECT 19.33 19.76 19.53 19.96 ;
        RECT 19.33 15.68 19.53 15.88 ;
        RECT 19.33 11.6 19.53 11.8 ;
        RECT 22.09 56.48 22.29 56.68 ;
        RECT 22.09 52.4 22.29 52.6 ;
        RECT 22.09 48.32 22.29 48.52 ;
        RECT 22.09 44.24 22.29 44.44 ;
        RECT 22.09 40.16 22.29 40.36 ;
        RECT 22.09 36.08 22.29 36.28 ;
        RECT 22.09 32 22.29 32.2 ;
        RECT 22.09 27.92 22.29 28.12 ;
        RECT 22.09 23.84 22.29 24.04 ;
        RECT 22.09 19.76 22.29 19.96 ;
        RECT 22.09 15.68 22.29 15.88 ;
        RECT 22.09 11.6 22.29 11.8 ;
        RECT 24.85 56.48 25.05 56.68 ;
        RECT 24.85 52.4 25.05 52.6 ;
        RECT 24.85 48.32 25.05 48.52 ;
        RECT 24.85 44.24 25.05 44.44 ;
        RECT 24.85 40.16 25.05 40.36 ;
        RECT 24.85 36.08 25.05 36.28 ;
        RECT 24.85 32 25.05 32.2 ;
        RECT 24.85 27.92 25.05 28.12 ;
        RECT 24.85 23.84 25.05 24.04 ;
        RECT 24.85 19.76 25.05 19.96 ;
        RECT 24.85 15.68 25.05 15.88 ;
        RECT 24.85 11.6 25.05 11.8 ;
        RECT 27.61 56.48 27.81 56.68 ;
        RECT 27.61 52.4 27.81 52.6 ;
        RECT 27.61 48.32 27.81 48.52 ;
        RECT 27.61 44.24 27.81 44.44 ;
        RECT 27.61 40.16 27.81 40.36 ;
        RECT 27.61 36.08 27.81 36.28 ;
        RECT 27.61 32 27.81 32.2 ;
        RECT 27.61 27.92 27.81 28.12 ;
        RECT 27.61 23.84 27.81 24.04 ;
        RECT 27.61 19.76 27.81 19.96 ;
        RECT 27.61 15.68 27.81 15.88 ;
        RECT 27.61 11.6 27.81 11.8 ;
        RECT 30.37 56.48 30.57 56.68 ;
        RECT 30.37 52.4 30.57 52.6 ;
        RECT 30.37 48.32 30.57 48.52 ;
        RECT 30.37 44.24 30.57 44.44 ;
        RECT 30.37 40.16 30.57 40.36 ;
        RECT 30.37 36.08 30.57 36.28 ;
        RECT 30.37 32 30.57 32.2 ;
        RECT 30.37 27.92 30.57 28.12 ;
        RECT 30.37 23.84 30.57 24.04 ;
        RECT 30.37 19.76 30.57 19.96 ;
        RECT 30.37 15.68 30.57 15.88 ;
        RECT 30.37 11.6 30.57 11.8 ;
        RECT 33.13 56.48 33.33 56.68 ;
        RECT 33.13 52.4 33.33 52.6 ;
        RECT 33.13 48.32 33.33 48.52 ;
        RECT 33.13 44.24 33.33 44.44 ;
        RECT 33.13 40.16 33.33 40.36 ;
        RECT 33.13 36.08 33.33 36.28 ;
        RECT 33.13 32 33.33 32.2 ;
        RECT 33.13 27.92 33.33 28.12 ;
        RECT 33.13 23.84 33.33 24.04 ;
        RECT 33.13 19.76 33.33 19.96 ;
        RECT 33.13 15.68 33.33 15.88 ;
        RECT 33.13 11.6 33.33 11.8 ;
        RECT 35.89 56.48 36.09 56.68 ;
        RECT 35.89 52.4 36.09 52.6 ;
        RECT 35.89 48.32 36.09 48.52 ;
        RECT 35.89 44.24 36.09 44.44 ;
        RECT 35.89 40.16 36.09 40.36 ;
        RECT 35.89 36.08 36.09 36.28 ;
        RECT 35.89 32 36.09 32.2 ;
        RECT 35.89 27.92 36.09 28.12 ;
        RECT 35.89 23.84 36.09 24.04 ;
        RECT 35.89 19.76 36.09 19.96 ;
        RECT 35.89 15.68 36.09 15.88 ;
        RECT 35.89 11.6 36.09 11.8 ;
        RECT 38.65 56.48 38.85 56.68 ;
        RECT 38.65 52.4 38.85 52.6 ;
        RECT 38.65 48.32 38.85 48.52 ;
        RECT 38.65 44.24 38.85 44.44 ;
        RECT 38.65 40.16 38.85 40.36 ;
        RECT 38.65 36.08 38.85 36.28 ;
        RECT 38.65 32 38.85 32.2 ;
        RECT 38.65 27.92 38.85 28.12 ;
        RECT 38.65 23.84 38.85 24.04 ;
        RECT 38.65 19.76 38.85 19.96 ;
        RECT 38.65 15.68 38.85 15.88 ;
        RECT 38.65 11.6 38.85 11.8 ;
        RECT 41.41 56.48 41.61 56.68 ;
        RECT 41.41 52.4 41.61 52.6 ;
        RECT 41.41 48.32 41.61 48.52 ;
        RECT 41.41 44.24 41.61 44.44 ;
        RECT 41.41 40.16 41.61 40.36 ;
        RECT 41.41 36.08 41.61 36.28 ;
        RECT 41.41 32 41.61 32.2 ;
        RECT 41.41 27.92 41.61 28.12 ;
        RECT 41.41 23.84 41.61 24.04 ;
        RECT 41.41 19.76 41.61 19.96 ;
        RECT 41.41 15.68 41.61 15.88 ;
        RECT 41.41 11.6 41.61 11.8 ;
        RECT 44.17 56.48 44.37 56.68 ;
        RECT 44.17 52.4 44.37 52.6 ;
        RECT 44.17 48.32 44.37 48.52 ;
        RECT 44.17 44.24 44.37 44.44 ;
        RECT 44.17 40.16 44.37 40.36 ;
        RECT 44.17 36.08 44.37 36.28 ;
        RECT 44.17 32 44.37 32.2 ;
        RECT 44.17 27.92 44.37 28.12 ;
        RECT 44.17 23.84 44.37 24.04 ;
        RECT 44.17 19.76 44.37 19.96 ;
        RECT 44.17 15.68 44.37 15.88 ;
        RECT 44.17 11.6 44.37 11.8 ;
        RECT 46.93 56.48 47.13 56.68 ;
        RECT 46.93 52.4 47.13 52.6 ;
        RECT 46.93 48.32 47.13 48.52 ;
        RECT 46.93 44.24 47.13 44.44 ;
        RECT 46.93 40.16 47.13 40.36 ;
        RECT 46.93 36.08 47.13 36.28 ;
        RECT 46.93 32 47.13 32.2 ;
        RECT 46.93 27.92 47.13 28.12 ;
        RECT 46.93 23.84 47.13 24.04 ;
        RECT 46.93 19.76 47.13 19.96 ;
        RECT 46.93 15.68 47.13 15.88 ;
        RECT 46.93 11.6 47.13 11.8 ;
        RECT 49.69 56.48 49.89 56.68 ;
        RECT 49.69 52.4 49.89 52.6 ;
        RECT 49.69 48.32 49.89 48.52 ;
        RECT 49.69 44.24 49.89 44.44 ;
        RECT 49.69 40.16 49.89 40.36 ;
        RECT 49.69 36.08 49.89 36.28 ;
        RECT 49.69 32 49.89 32.2 ;
        RECT 49.69 27.92 49.89 28.12 ;
        RECT 49.69 23.84 49.89 24.04 ;
        RECT 49.69 19.76 49.89 19.96 ;
        RECT 49.69 15.68 49.89 15.88 ;
        RECT 49.69 11.6 49.89 11.8 ;
        RECT 52.45 56.48 52.65 56.68 ;
        RECT 52.45 52.4 52.65 52.6 ;
        RECT 52.45 48.32 52.65 48.52 ;
        RECT 52.45 44.24 52.65 44.44 ;
        RECT 52.45 40.16 52.65 40.36 ;
        RECT 52.45 36.08 52.65 36.28 ;
        RECT 52.45 32 52.65 32.2 ;
        RECT 52.45 27.92 52.65 28.12 ;
        RECT 52.45 23.84 52.65 24.04 ;
        RECT 52.45 19.76 52.65 19.96 ;
        RECT 52.45 15.68 52.65 15.88 ;
        RECT 52.45 11.6 52.65 11.8 ;
        RECT 55.21 56.48 55.41 56.68 ;
        RECT 55.21 52.4 55.41 52.6 ;
        RECT 55.21 48.32 55.41 48.52 ;
        RECT 55.21 44.24 55.41 44.44 ;
        RECT 55.21 40.16 55.41 40.36 ;
        RECT 55.21 36.08 55.41 36.28 ;
        RECT 55.21 32 55.41 32.2 ;
        RECT 55.21 27.92 55.41 28.12 ;
        RECT 55.21 23.84 55.41 24.04 ;
        RECT 55.21 19.76 55.41 19.96 ;
        RECT 55.21 15.68 55.41 15.88 ;
        RECT 55.21 11.6 55.41 11.8 ;
        RECT 57.97 56.48 58.17 56.68 ;
        RECT 57.97 52.4 58.17 52.6 ;
        RECT 57.97 48.32 58.17 48.52 ;
        RECT 57.97 44.24 58.17 44.44 ;
        RECT 57.97 40.16 58.17 40.36 ;
        RECT 57.97 36.08 58.17 36.28 ;
        RECT 57.97 32 58.17 32.2 ;
        RECT 57.97 27.92 58.17 28.12 ;
        RECT 57.97 23.84 58.17 24.04 ;
        RECT 57.97 19.76 58.17 19.96 ;
        RECT 57.97 15.68 58.17 15.88 ;
        RECT 57.97 11.6 58.17 11.8 ;
        RECT 60.73 56.48 60.93 56.68 ;
        RECT 60.73 52.4 60.93 52.6 ;
        RECT 60.73 48.32 60.93 48.52 ;
        RECT 60.73 44.24 60.93 44.44 ;
        RECT 60.73 40.16 60.93 40.36 ;
        RECT 60.73 36.08 60.93 36.28 ;
        RECT 60.73 32 60.93 32.2 ;
        RECT 60.73 27.92 60.93 28.12 ;
        RECT 60.73 23.84 60.93 24.04 ;
        RECT 60.73 19.76 60.93 19.96 ;
        RECT 60.73 15.68 60.93 15.88 ;
        RECT 60.73 11.6 60.93 11.8 ;
        RECT 63.49 56.48 63.69 56.68 ;
        RECT 63.49 52.4 63.69 52.6 ;
        RECT 63.49 48.32 63.69 48.52 ;
        RECT 63.49 44.24 63.69 44.44 ;
        RECT 63.49 40.16 63.69 40.36 ;
        RECT 63.49 36.08 63.69 36.28 ;
        RECT 63.49 32 63.69 32.2 ;
        RECT 63.49 27.92 63.69 28.12 ;
        RECT 63.49 23.84 63.69 24.04 ;
        RECT 63.49 19.76 63.69 19.96 ;
        RECT 63.49 15.68 63.69 15.88 ;
        RECT 63.49 11.6 63.69 11.8 ;
        RECT 66.25 56.48 66.45 56.68 ;
        RECT 66.25 52.4 66.45 52.6 ;
        RECT 66.25 48.32 66.45 48.52 ;
        RECT 66.25 44.24 66.45 44.44 ;
        RECT 66.25 40.16 66.45 40.36 ;
        RECT 66.25 36.08 66.45 36.28 ;
        RECT 66.25 32 66.45 32.2 ;
        RECT 66.25 27.92 66.45 28.12 ;
        RECT 66.25 23.84 66.45 24.04 ;
        RECT 66.25 19.76 66.45 19.96 ;
        RECT 66.25 15.68 66.45 15.88 ;
        RECT 66.25 11.6 66.45 11.8 ;
        RECT 69.01 56.48 69.21 56.68 ;
        RECT 69.01 52.4 69.21 52.6 ;
        RECT 69.01 48.32 69.21 48.52 ;
        RECT 69.01 44.24 69.21 44.44 ;
        RECT 69.01 40.16 69.21 40.36 ;
        RECT 69.01 36.08 69.21 36.28 ;
        RECT 69.01 32 69.21 32.2 ;
        RECT 69.01 27.92 69.21 28.12 ;
        RECT 69.01 23.84 69.21 24.04 ;
        RECT 69.01 19.76 69.21 19.96 ;
        RECT 69.01 15.68 69.21 15.88 ;
        RECT 69.01 11.6 69.21 11.8 ;
        RECT 71.77 56.48 71.97 56.68 ;
        RECT 71.77 52.4 71.97 52.6 ;
        RECT 71.77 48.32 71.97 48.52 ;
        RECT 71.77 44.24 71.97 44.44 ;
        RECT 71.77 40.16 71.97 40.36 ;
        RECT 71.77 36.08 71.97 36.28 ;
        RECT 71.77 32 71.97 32.2 ;
        RECT 71.77 27.92 71.97 28.12 ;
        RECT 71.77 23.84 71.97 24.04 ;
        RECT 71.77 19.76 71.97 19.96 ;
        RECT 71.77 15.68 71.97 15.88 ;
        RECT 71.77 11.6 71.97 11.8 ;
        RECT 74.53 56.48 74.73 56.68 ;
        RECT 74.53 52.4 74.73 52.6 ;
        RECT 74.53 48.32 74.73 48.52 ;
        RECT 74.53 44.24 74.73 44.44 ;
        RECT 74.53 40.16 74.73 40.36 ;
        RECT 74.53 36.08 74.73 36.28 ;
        RECT 74.53 32 74.73 32.2 ;
        RECT 74.53 27.92 74.73 28.12 ;
        RECT 74.53 23.84 74.73 24.04 ;
        RECT 74.53 19.76 74.73 19.96 ;
        RECT 74.53 15.68 74.73 15.88 ;
        RECT 74.53 11.6 74.73 11.8 ;
        RECT 77.29 56.48 77.49 56.68 ;
        RECT 77.29 52.4 77.49 52.6 ;
        RECT 77.29 48.32 77.49 48.52 ;
        RECT 77.29 44.24 77.49 44.44 ;
        RECT 77.29 40.16 77.49 40.36 ;
        RECT 77.29 36.08 77.49 36.28 ;
        RECT 77.29 32 77.49 32.2 ;
        RECT 77.29 27.92 77.49 28.12 ;
        RECT 77.29 23.84 77.49 24.04 ;
        RECT 77.29 19.76 77.49 19.96 ;
        RECT 77.29 15.68 77.49 15.88 ;
        RECT 77.29 11.6 77.49 11.8 ;
        RECT 80.05 56.48 80.25 56.68 ;
        RECT 80.05 52.4 80.25 52.6 ;
        RECT 80.05 48.32 80.25 48.52 ;
        RECT 80.05 44.24 80.25 44.44 ;
        RECT 80.05 40.16 80.25 40.36 ;
        RECT 80.05 36.08 80.25 36.28 ;
        RECT 80.05 32 80.25 32.2 ;
        RECT 80.05 27.92 80.25 28.12 ;
        RECT 80.05 23.84 80.25 24.04 ;
        RECT 80.05 19.76 80.25 19.96 ;
        RECT 80.05 15.68 80.25 15.88 ;
        RECT 80.05 11.6 80.25 11.8 ;
        RECT 82.81 56.48 83.01 56.68 ;
        RECT 82.81 52.4 83.01 52.6 ;
        RECT 82.81 48.32 83.01 48.52 ;
        RECT 82.81 44.24 83.01 44.44 ;
        RECT 82.81 40.16 83.01 40.36 ;
        RECT 82.81 36.08 83.01 36.28 ;
        RECT 82.81 32 83.01 32.2 ;
        RECT 82.81 27.92 83.01 28.12 ;
        RECT 82.81 23.84 83.01 24.04 ;
        RECT 82.81 19.76 83.01 19.96 ;
        RECT 82.81 15.68 83.01 15.88 ;
        RECT 82.81 11.6 83.01 11.8 ;
        RECT 85.57 56.48 85.77 56.68 ;
        RECT 85.57 52.4 85.77 52.6 ;
        RECT 85.57 48.32 85.77 48.52 ;
        RECT 85.57 44.24 85.77 44.44 ;
        RECT 85.57 40.16 85.77 40.36 ;
        RECT 85.57 36.08 85.77 36.28 ;
        RECT 85.57 32 85.77 32.2 ;
        RECT 85.57 27.92 85.77 28.12 ;
        RECT 85.57 23.84 85.77 24.04 ;
        RECT 85.57 19.76 85.77 19.96 ;
        RECT 85.57 15.68 85.77 15.88 ;
        RECT 85.57 11.6 85.77 11.8 ;
        RECT 88.33 56.48 88.53 56.68 ;
        RECT 88.33 52.4 88.53 52.6 ;
        RECT 88.33 48.32 88.53 48.52 ;
        RECT 88.33 44.24 88.53 44.44 ;
        RECT 88.33 40.16 88.53 40.36 ;
        RECT 88.33 36.08 88.53 36.28 ;
        RECT 88.33 32 88.53 32.2 ;
        RECT 88.33 27.92 88.53 28.12 ;
        RECT 88.33 23.84 88.53 24.04 ;
        RECT 88.33 19.76 88.53 19.96 ;
        RECT 88.33 15.68 88.53 15.88 ;
        RECT 88.33 11.6 88.53 11.8 ;
        RECT 91.09 56.48 91.29 56.68 ;
        RECT 91.09 52.4 91.29 52.6 ;
        RECT 91.09 48.32 91.29 48.52 ;
        RECT 91.09 44.24 91.29 44.44 ;
        RECT 91.09 40.16 91.29 40.36 ;
        RECT 91.09 36.08 91.29 36.28 ;
        RECT 91.09 32 91.29 32.2 ;
        RECT 91.09 27.92 91.29 28.12 ;
        RECT 91.09 23.84 91.29 24.04 ;
        RECT 91.09 19.76 91.29 19.96 ;
        RECT 91.09 15.68 91.29 15.88 ;
        RECT 91.09 11.6 91.29 11.8 ;
        RECT 93.85 56.48 94.05 56.68 ;
        RECT 93.85 52.4 94.05 52.6 ;
        RECT 93.85 48.32 94.05 48.52 ;
        RECT 93.85 44.24 94.05 44.44 ;
        RECT 93.85 40.16 94.05 40.36 ;
        RECT 93.85 36.08 94.05 36.28 ;
        RECT 93.85 32 94.05 32.2 ;
        RECT 93.85 27.92 94.05 28.12 ;
        RECT 93.85 23.84 94.05 24.04 ;
        RECT 93.85 19.76 94.05 19.96 ;
        RECT 93.85 15.68 94.05 15.88 ;
        RECT 93.85 11.6 94.05 11.8 ;
        RECT 96.61 56.48 96.81 56.68 ;
        RECT 96.61 52.4 96.81 52.6 ;
        RECT 96.61 48.32 96.81 48.52 ;
        RECT 96.61 44.24 96.81 44.44 ;
        RECT 96.61 40.16 96.81 40.36 ;
        RECT 96.61 36.08 96.81 36.28 ;
        RECT 96.61 32 96.81 32.2 ;
        RECT 96.61 27.92 96.81 28.12 ;
        RECT 96.61 23.84 96.81 24.04 ;
        RECT 96.61 19.76 96.81 19.96 ;
        RECT 96.61 15.68 96.81 15.88 ;
        RECT 96.61 11.6 96.81 11.8 ;
        RECT 99.37 56.48 99.57 56.68 ;
        RECT 99.37 52.4 99.57 52.6 ;
        RECT 99.37 48.32 99.57 48.52 ;
        RECT 99.37 44.24 99.57 44.44 ;
        RECT 99.37 40.16 99.57 40.36 ;
        RECT 99.37 36.08 99.57 36.28 ;
        RECT 99.37 32 99.57 32.2 ;
        RECT 99.37 27.92 99.57 28.12 ;
        RECT 99.37 23.84 99.57 24.04 ;
        RECT 99.37 19.76 99.57 19.96 ;
        RECT 99.37 15.68 99.57 15.88 ;
        RECT 99.37 11.6 99.57 11.8 ;
        RECT 102.13 56.48 102.33 56.68 ;
        RECT 102.13 52.4 102.33 52.6 ;
        RECT 102.13 48.32 102.33 48.52 ;
        RECT 102.13 44.24 102.33 44.44 ;
        RECT 102.13 40.16 102.33 40.36 ;
        RECT 102.13 36.08 102.33 36.28 ;
        RECT 102.13 32 102.33 32.2 ;
        RECT 102.13 27.92 102.33 28.12 ;
        RECT 102.13 23.84 102.33 24.04 ;
        RECT 102.13 19.76 102.33 19.96 ;
        RECT 102.13 15.68 102.33 15.88 ;
        RECT 102.13 11.6 102.33 11.8 ;
        RECT 104.89 56.48 105.09 56.68 ;
        RECT 104.89 52.4 105.09 52.6 ;
        RECT 104.89 48.32 105.09 48.52 ;
        RECT 104.89 44.24 105.09 44.44 ;
        RECT 104.89 40.16 105.09 40.36 ;
        RECT 104.89 36.08 105.09 36.28 ;
        RECT 104.89 32 105.09 32.2 ;
        RECT 104.89 27.92 105.09 28.12 ;
        RECT 104.89 23.84 105.09 24.04 ;
        RECT 104.89 19.76 105.09 19.96 ;
        RECT 104.89 15.68 105.09 15.88 ;
        RECT 104.89 11.6 105.09 11.8 ;
        RECT 107.65 56.48 107.85 56.68 ;
        RECT 107.65 52.4 107.85 52.6 ;
        RECT 107.65 48.32 107.85 48.52 ;
        RECT 107.65 44.24 107.85 44.44 ;
        RECT 107.65 40.16 107.85 40.36 ;
        RECT 107.65 36.08 107.85 36.28 ;
        RECT 107.65 32 107.85 32.2 ;
        RECT 107.65 27.92 107.85 28.12 ;
        RECT 107.65 23.84 107.85 24.04 ;
        RECT 107.65 19.76 107.85 19.96 ;
        RECT 107.65 15.68 107.85 15.88 ;
        RECT 107.65 11.6 107.85 11.8 ;
        RECT 110.41 56.48 110.61 56.68 ;
        RECT 110.41 52.4 110.61 52.6 ;
        RECT 110.41 48.32 110.61 48.52 ;
        RECT 110.41 44.24 110.61 44.44 ;
        RECT 110.41 40.16 110.61 40.36 ;
        RECT 110.41 36.08 110.61 36.28 ;
        RECT 110.41 32 110.61 32.2 ;
        RECT 110.41 27.92 110.61 28.12 ;
        RECT 110.41 23.84 110.61 24.04 ;
        RECT 110.41 19.76 110.61 19.96 ;
        RECT 110.41 15.68 110.61 15.88 ;
        RECT 110.41 11.6 110.61 11.8 ;
        RECT 113.17 56.48 113.37 56.68 ;
        RECT 113.17 52.4 113.37 52.6 ;
        RECT 113.17 48.32 113.37 48.52 ;
        RECT 113.17 44.24 113.37 44.44 ;
        RECT 113.17 40.16 113.37 40.36 ;
        RECT 113.17 36.08 113.37 36.28 ;
        RECT 113.17 32 113.37 32.2 ;
        RECT 113.17 27.92 113.37 28.12 ;
        RECT 113.17 23.84 113.37 24.04 ;
        RECT 113.17 19.76 113.37 19.96 ;
        RECT 113.17 15.68 113.37 15.88 ;
        RECT 113.17 11.6 113.37 11.8 ;
        RECT 115.93 56.48 116.13 56.68 ;
        RECT 115.93 52.4 116.13 52.6 ;
        RECT 115.93 48.32 116.13 48.52 ;
        RECT 115.93 44.24 116.13 44.44 ;
        RECT 115.93 40.16 116.13 40.36 ;
        RECT 115.93 36.08 116.13 36.28 ;
        RECT 115.93 32 116.13 32.2 ;
        RECT 115.93 27.92 116.13 28.12 ;
        RECT 115.93 23.84 116.13 24.04 ;
        RECT 115.93 19.76 116.13 19.96 ;
        RECT 115.93 15.68 116.13 15.88 ;
        RECT 115.93 11.6 116.13 11.8 ;
        RECT 118.69 56.48 118.89 56.68 ;
        RECT 118.69 52.4 118.89 52.6 ;
        RECT 118.69 48.32 118.89 48.52 ;
        RECT 118.69 44.24 118.89 44.44 ;
        RECT 118.69 40.16 118.89 40.36 ;
        RECT 118.69 36.08 118.89 36.28 ;
        RECT 118.69 32 118.89 32.2 ;
        RECT 118.69 27.92 118.89 28.12 ;
        RECT 118.69 23.84 118.89 24.04 ;
        RECT 118.69 19.76 118.89 19.96 ;
        RECT 118.69 15.68 118.89 15.88 ;
        RECT 118.69 11.6 118.89 11.8 ;
        RECT 121.45 56.48 121.65 56.68 ;
        RECT 121.45 52.4 121.65 52.6 ;
        RECT 121.45 48.32 121.65 48.52 ;
        RECT 121.45 44.24 121.65 44.44 ;
        RECT 121.45 40.16 121.65 40.36 ;
        RECT 121.45 36.08 121.65 36.28 ;
        RECT 121.45 32 121.65 32.2 ;
        RECT 121.45 27.92 121.65 28.12 ;
        RECT 121.45 23.84 121.65 24.04 ;
        RECT 121.45 19.76 121.65 19.96 ;
        RECT 121.45 15.68 121.65 15.88 ;
        RECT 121.45 11.6 121.65 11.8 ;
        RECT 124.21 56.48 124.41 56.68 ;
        RECT 124.21 52.4 124.41 52.6 ;
        RECT 124.21 48.32 124.41 48.52 ;
        RECT 124.21 44.24 124.41 44.44 ;
        RECT 124.21 40.16 124.41 40.36 ;
        RECT 124.21 36.08 124.41 36.28 ;
        RECT 124.21 32 124.41 32.2 ;
        RECT 124.21 27.92 124.41 28.12 ;
        RECT 124.21 23.84 124.41 24.04 ;
        RECT 124.21 19.76 124.41 19.96 ;
        RECT 124.21 15.68 124.41 15.88 ;
        RECT 124.21 11.6 124.41 11.8 ;
        RECT 126.97 56.48 127.17 56.68 ;
        RECT 126.97 52.4 127.17 52.6 ;
        RECT 126.97 48.32 127.17 48.52 ;
        RECT 126.97 44.24 127.17 44.44 ;
        RECT 126.97 40.16 127.17 40.36 ;
        RECT 126.97 36.08 127.17 36.28 ;
        RECT 126.97 32 127.17 32.2 ;
        RECT 126.97 27.92 127.17 28.12 ;
        RECT 126.97 23.84 127.17 24.04 ;
        RECT 126.97 19.76 127.17 19.96 ;
        RECT 126.97 15.68 127.17 15.88 ;
        RECT 126.97 11.6 127.17 11.8 ;
        RECT 129.73 56.48 129.93 56.68 ;
        RECT 129.73 52.4 129.93 52.6 ;
        RECT 129.73 48.32 129.93 48.52 ;
        RECT 129.73 44.24 129.93 44.44 ;
        RECT 129.73 40.16 129.93 40.36 ;
        RECT 129.73 36.08 129.93 36.28 ;
        RECT 129.73 32 129.93 32.2 ;
        RECT 129.73 27.92 129.93 28.12 ;
        RECT 129.73 23.84 129.93 24.04 ;
        RECT 129.73 19.76 129.93 19.96 ;
        RECT 129.73 15.68 129.93 15.88 ;
        RECT 129.73 11.6 129.93 11.8 ;
        RECT 132.49 56.48 132.69 56.68 ;
        RECT 132.49 52.4 132.69 52.6 ;
        RECT 132.49 48.32 132.69 48.52 ;
        RECT 132.49 44.24 132.69 44.44 ;
        RECT 132.49 40.16 132.69 40.36 ;
        RECT 132.49 36.08 132.69 36.28 ;
        RECT 132.49 32 132.69 32.2 ;
        RECT 132.49 27.92 132.69 28.12 ;
        RECT 132.49 23.84 132.69 24.04 ;
        RECT 132.49 19.76 132.69 19.96 ;
        RECT 132.49 15.68 132.69 15.88 ;
        RECT 132.49 11.6 132.69 11.8 ;
        RECT 135.25 56.48 135.45 56.68 ;
        RECT 135.25 52.4 135.45 52.6 ;
        RECT 135.25 48.32 135.45 48.52 ;
        RECT 135.25 44.24 135.45 44.44 ;
        RECT 135.25 40.16 135.45 40.36 ;
        RECT 135.25 36.08 135.45 36.28 ;
        RECT 135.25 32 135.45 32.2 ;
        RECT 135.25 27.92 135.45 28.12 ;
        RECT 135.25 23.84 135.45 24.04 ;
        RECT 135.25 19.76 135.45 19.96 ;
        RECT 135.25 15.68 135.45 15.88 ;
        RECT 135.25 11.6 135.45 11.8 ;
        RECT 138.01 56.48 138.21 56.68 ;
        RECT 138.01 52.4 138.21 52.6 ;
        RECT 138.01 48.32 138.21 48.52 ;
        RECT 138.01 44.24 138.21 44.44 ;
        RECT 138.01 40.16 138.21 40.36 ;
        RECT 138.01 36.08 138.21 36.28 ;
        RECT 138.01 32 138.21 32.2 ;
        RECT 138.01 27.92 138.21 28.12 ;
        RECT 138.01 23.84 138.21 24.04 ;
        RECT 138.01 19.76 138.21 19.96 ;
        RECT 138.01 15.68 138.21 15.88 ;
        RECT 138.01 11.6 138.21 11.8 ;
        RECT 140.77 56.48 140.97 56.68 ;
        RECT 140.77 52.4 140.97 52.6 ;
        RECT 140.77 48.32 140.97 48.52 ;
        RECT 140.77 44.24 140.97 44.44 ;
        RECT 140.77 40.16 140.97 40.36 ;
        RECT 140.77 36.08 140.97 36.28 ;
        RECT 140.77 32 140.97 32.2 ;
        RECT 140.77 27.92 140.97 28.12 ;
        RECT 140.77 23.84 140.97 24.04 ;
        RECT 140.77 19.76 140.97 19.96 ;
        RECT 140.77 15.68 140.97 15.88 ;
        RECT 140.77 11.6 140.97 11.8 ;
        RECT 143.53 56.48 143.73 56.68 ;
        RECT 143.53 52.4 143.73 52.6 ;
        RECT 143.53 48.32 143.73 48.52 ;
        RECT 143.53 44.24 143.73 44.44 ;
        RECT 143.53 40.16 143.73 40.36 ;
        RECT 143.53 36.08 143.73 36.28 ;
        RECT 143.53 32 143.73 32.2 ;
        RECT 143.53 27.92 143.73 28.12 ;
        RECT 143.53 23.84 143.73 24.04 ;
        RECT 143.53 19.76 143.73 19.96 ;
        RECT 143.53 15.68 143.73 15.88 ;
        RECT 143.53 11.6 143.73 11.8 ;
        RECT 146.29 56.48 146.49 56.68 ;
        RECT 146.29 52.4 146.49 52.6 ;
        RECT 146.29 48.32 146.49 48.52 ;
        RECT 146.29 44.24 146.49 44.44 ;
        RECT 146.29 40.16 146.49 40.36 ;
        RECT 146.29 36.08 146.49 36.28 ;
        RECT 146.29 32 146.49 32.2 ;
        RECT 146.29 27.92 146.49 28.12 ;
        RECT 146.29 23.84 146.49 24.04 ;
        RECT 146.29 19.76 146.49 19.96 ;
        RECT 146.29 15.68 146.49 15.88 ;
        RECT 146.29 11.6 146.49 11.8 ;
        RECT 149.05 56.48 149.25 56.68 ;
        RECT 149.05 52.4 149.25 52.6 ;
        RECT 149.05 48.32 149.25 48.52 ;
        RECT 149.05 44.24 149.25 44.44 ;
        RECT 149.05 40.16 149.25 40.36 ;
        RECT 149.05 36.08 149.25 36.28 ;
        RECT 149.05 32 149.25 32.2 ;
        RECT 149.05 27.92 149.25 28.12 ;
        RECT 149.05 23.84 149.25 24.04 ;
        RECT 149.05 19.76 149.25 19.96 ;
        RECT 149.05 15.68 149.25 15.88 ;
        RECT 149.05 11.6 149.25 11.8 ;
        RECT 151.81 56.48 152.01 56.68 ;
        RECT 151.81 52.4 152.01 52.6 ;
        RECT 151.81 48.32 152.01 48.52 ;
        RECT 151.81 44.24 152.01 44.44 ;
        RECT 151.81 40.16 152.01 40.36 ;
        RECT 151.81 36.08 152.01 36.28 ;
        RECT 151.81 32 152.01 32.2 ;
        RECT 151.81 27.92 152.01 28.12 ;
        RECT 151.81 23.84 152.01 24.04 ;
        RECT 151.81 19.76 152.01 19.96 ;
        RECT 151.81 15.68 152.01 15.88 ;
        RECT 151.81 11.6 152.01 11.8 ;
        RECT 154.57 56.48 154.77 56.68 ;
        RECT 154.57 52.4 154.77 52.6 ;
        RECT 154.57 48.32 154.77 48.52 ;
        RECT 154.57 44.24 154.77 44.44 ;
        RECT 154.57 40.16 154.77 40.36 ;
        RECT 154.57 36.08 154.77 36.28 ;
        RECT 154.57 32 154.77 32.2 ;
        RECT 154.57 27.92 154.77 28.12 ;
        RECT 154.57 23.84 154.77 24.04 ;
        RECT 154.57 19.76 154.77 19.96 ;
        RECT 154.57 15.68 154.77 15.88 ;
        RECT 154.57 11.6 154.77 11.8 ;
        RECT 157.33 56.48 157.53 56.68 ;
        RECT 157.33 52.4 157.53 52.6 ;
        RECT 157.33 48.32 157.53 48.52 ;
        RECT 157.33 44.24 157.53 44.44 ;
        RECT 157.33 40.16 157.53 40.36 ;
        RECT 157.33 36.08 157.53 36.28 ;
        RECT 157.33 32 157.53 32.2 ;
        RECT 157.33 27.92 157.53 28.12 ;
        RECT 157.33 23.84 157.53 24.04 ;
        RECT 157.33 19.76 157.53 19.96 ;
        RECT 157.33 15.68 157.53 15.88 ;
        RECT 157.33 11.6 157.53 11.8 ;
        RECT 160.09 56.48 160.29 56.68 ;
        RECT 160.09 52.4 160.29 52.6 ;
        RECT 160.09 48.32 160.29 48.52 ;
        RECT 160.09 44.24 160.29 44.44 ;
        RECT 160.09 40.16 160.29 40.36 ;
        RECT 160.09 36.08 160.29 36.28 ;
        RECT 160.09 32 160.29 32.2 ;
        RECT 160.09 27.92 160.29 28.12 ;
        RECT 160.09 23.84 160.29 24.04 ;
        RECT 160.09 19.76 160.29 19.96 ;
        RECT 160.09 15.68 160.29 15.88 ;
        RECT 160.09 11.6 160.29 11.8 ;
        RECT 162.85 56.48 163.05 56.68 ;
        RECT 162.85 52.4 163.05 52.6 ;
        RECT 162.85 48.32 163.05 48.52 ;
        RECT 162.85 44.24 163.05 44.44 ;
        RECT 162.85 40.16 163.05 40.36 ;
        RECT 162.85 36.08 163.05 36.28 ;
        RECT 162.85 32 163.05 32.2 ;
        RECT 162.85 27.92 163.05 28.12 ;
        RECT 162.85 23.84 163.05 24.04 ;
        RECT 162.85 19.76 163.05 19.96 ;
        RECT 162.85 15.68 163.05 15.88 ;
        RECT 162.85 11.6 163.05 11.8 ;
        RECT 165.61 56.48 165.81 56.68 ;
        RECT 165.61 52.4 165.81 52.6 ;
        RECT 165.61 48.32 165.81 48.52 ;
        RECT 165.61 44.24 165.81 44.44 ;
        RECT 165.61 40.16 165.81 40.36 ;
        RECT 165.61 36.08 165.81 36.28 ;
        RECT 165.61 32 165.81 32.2 ;
        RECT 165.61 27.92 165.81 28.12 ;
        RECT 165.61 23.84 165.81 24.04 ;
        RECT 165.61 19.76 165.81 19.96 ;
        RECT 165.61 15.68 165.81 15.88 ;
        RECT 165.61 11.6 165.81 11.8 ;
        RECT 168.37 56.48 168.57 56.68 ;
        RECT 168.37 52.4 168.57 52.6 ;
        RECT 168.37 48.32 168.57 48.52 ;
        RECT 168.37 44.24 168.57 44.44 ;
        RECT 168.37 40.16 168.57 40.36 ;
        RECT 168.37 36.08 168.57 36.28 ;
        RECT 168.37 32 168.57 32.2 ;
        RECT 168.37 27.92 168.57 28.12 ;
        RECT 168.37 23.84 168.57 24.04 ;
        RECT 168.37 19.76 168.57 19.96 ;
        RECT 168.37 15.68 168.57 15.88 ;
        RECT 168.37 11.6 168.57 11.8 ;
        RECT 171.13 56.48 171.33 56.68 ;
        RECT 171.13 52.4 171.33 52.6 ;
        RECT 171.13 48.32 171.33 48.52 ;
        RECT 171.13 44.24 171.33 44.44 ;
        RECT 171.13 40.16 171.33 40.36 ;
        RECT 171.13 36.08 171.33 36.28 ;
        RECT 171.13 32 171.33 32.2 ;
        RECT 171.13 27.92 171.33 28.12 ;
        RECT 171.13 23.84 171.33 24.04 ;
        RECT 171.13 19.76 171.33 19.96 ;
        RECT 171.13 15.68 171.33 15.88 ;
        RECT 171.13 11.6 171.33 11.8 ;
        RECT 173.89 56.48 174.09 56.68 ;
        RECT 173.89 52.4 174.09 52.6 ;
        RECT 173.89 48.32 174.09 48.52 ;
        RECT 173.89 44.24 174.09 44.44 ;
        RECT 173.89 40.16 174.09 40.36 ;
        RECT 173.89 36.08 174.09 36.28 ;
        RECT 173.89 32 174.09 32.2 ;
        RECT 173.89 27.92 174.09 28.12 ;
        RECT 173.89 23.84 174.09 24.04 ;
        RECT 173.89 19.76 174.09 19.96 ;
        RECT 173.89 15.68 174.09 15.88 ;
        RECT 173.89 11.6 174.09 11.8 ;
        RECT 176.65 56.48 176.85 56.68 ;
        RECT 176.65 52.4 176.85 52.6 ;
        RECT 176.65 48.32 176.85 48.52 ;
        RECT 176.65 44.24 176.85 44.44 ;
        RECT 176.65 40.16 176.85 40.36 ;
        RECT 176.65 36.08 176.85 36.28 ;
        RECT 176.65 32 176.85 32.2 ;
        RECT 176.65 27.92 176.85 28.12 ;
        RECT 176.65 23.84 176.85 24.04 ;
        RECT 176.65 19.76 176.85 19.96 ;
        RECT 176.65 15.68 176.85 15.88 ;
        RECT 176.65 11.6 176.85 11.8 ;
        RECT 179.41 56.48 179.61 56.68 ;
        RECT 179.41 52.4 179.61 52.6 ;
        RECT 179.41 48.32 179.61 48.52 ;
        RECT 179.41 44.24 179.61 44.44 ;
        RECT 179.41 40.16 179.61 40.36 ;
        RECT 179.41 36.08 179.61 36.28 ;
        RECT 179.41 32 179.61 32.2 ;
        RECT 179.41 27.92 179.61 28.12 ;
        RECT 179.41 23.84 179.61 24.04 ;
        RECT 179.41 19.76 179.61 19.96 ;
        RECT 179.41 15.68 179.61 15.88 ;
        RECT 179.41 11.6 179.61 11.8 ;
        RECT 182.17 56.48 182.37 56.68 ;
        RECT 182.17 52.4 182.37 52.6 ;
        RECT 182.17 48.32 182.37 48.52 ;
        RECT 182.17 44.24 182.37 44.44 ;
        RECT 182.17 40.16 182.37 40.36 ;
        RECT 182.17 36.08 182.37 36.28 ;
        RECT 182.17 32 182.37 32.2 ;
        RECT 182.17 27.92 182.37 28.12 ;
        RECT 182.17 23.84 182.37 24.04 ;
        RECT 182.17 19.76 182.37 19.96 ;
        RECT 182.17 15.68 182.37 15.88 ;
        RECT 182.17 11.6 182.37 11.8 ;
        RECT 184.93 56.48 185.13 56.68 ;
        RECT 184.93 52.4 185.13 52.6 ;
        RECT 184.93 48.32 185.13 48.52 ;
        RECT 184.93 44.24 185.13 44.44 ;
        RECT 184.93 40.16 185.13 40.36 ;
        RECT 184.93 36.08 185.13 36.28 ;
        RECT 184.93 32 185.13 32.2 ;
        RECT 184.93 27.92 185.13 28.12 ;
        RECT 184.93 23.84 185.13 24.04 ;
        RECT 184.93 19.76 185.13 19.96 ;
        RECT 184.93 15.68 185.13 15.88 ;
        RECT 184.93 11.6 185.13 11.8 ;
        RECT 187.69 56.48 187.89 56.68 ;
        RECT 187.69 52.4 187.89 52.6 ;
        RECT 187.69 48.32 187.89 48.52 ;
        RECT 187.69 44.24 187.89 44.44 ;
        RECT 187.69 40.16 187.89 40.36 ;
        RECT 187.69 36.08 187.89 36.28 ;
        RECT 187.69 32 187.89 32.2 ;
        RECT 187.69 27.92 187.89 28.12 ;
        RECT 187.69 23.84 187.89 24.04 ;
        RECT 187.69 19.76 187.89 19.96 ;
        RECT 187.69 15.68 187.89 15.88 ;
        RECT 187.69 11.6 187.89 11.8 ;
    END
  END VSS
  OBS
    LAYER mcon ;
      RECT 184.025 21.305 184.195 21.475 ;
      RECT 181.715 21.985 181.885 22.155 ;
      RECT 181.28 21.645 181.45 21.815 ;
      RECT 181.265 24.705 181.435 24.875 ;
      RECT 179.71 21.645 179.88 21.815 ;
      RECT 179.195 21.985 179.365 22.155 ;
      RECT 178.43 22.665 178.6 22.835 ;
      RECT 178.005 21.985 178.175 22.155 ;
      RECT 177.61 21.645 177.78 21.815 ;
      RECT 177.125 16.885 177.295 17.055 ;
      RECT 177.125 21.985 177.295 22.155 ;
      RECT 176.205 15.865 176.375 16.035 ;
      RECT 173.905 20.285 174.075 20.455 ;
      RECT 173.895 16.545 174.065 16.715 ;
      RECT 173.46 16.205 173.63 16.375 ;
      RECT 172.985 22.665 173.155 22.835 ;
      RECT 172.525 19.945 172.695 20.115 ;
      RECT 171.89 16.205 172.06 16.375 ;
      RECT 171.605 24.705 171.775 24.875 ;
      RECT 171.375 16.545 171.545 16.715 ;
      RECT 171.145 21.645 171.315 21.815 ;
      RECT 171.145 24.025 171.315 24.195 ;
      RECT 170.64 16.885 170.81 17.055 ;
      RECT 170.225 24.705 170.395 24.875 ;
      RECT 170.215 19.605 170.385 19.775 ;
      RECT 170.185 16.545 170.355 16.715 ;
      RECT 169.79 16.205 169.96 16.375 ;
      RECT 169.78 19.945 169.95 20.115 ;
      RECT 169.765 13.825 169.935 13.995 ;
      RECT 169.305 13.485 169.475 13.655 ;
      RECT 169.305 16.885 169.475 17.055 ;
      RECT 169.305 21.305 169.475 21.475 ;
      RECT 169.305 23.005 169.475 23.175 ;
      RECT 169.305 24.365 169.475 24.535 ;
      RECT 168.615 13.825 168.785 13.995 ;
      RECT 168.21 19.945 168.38 20.115 ;
      RECT 167.925 14.845 168.095 15.015 ;
      RECT 167.695 19.605 167.865 19.775 ;
      RECT 166.995 21.985 167.165 22.155 ;
      RECT 166.93 18.925 167.1 19.095 ;
      RECT 166.56 21.645 166.73 21.815 ;
      RECT 166.505 19.605 166.675 19.775 ;
      RECT 166.11 19.945 166.28 20.115 ;
      RECT 165.625 19.265 165.795 19.435 ;
      RECT 165.165 18.925 165.335 19.095 ;
      RECT 164.99 21.645 165.16 21.815 ;
      RECT 164.475 21.985 164.645 22.155 ;
      RECT 164.245 11.445 164.415 11.615 ;
      RECT 163.71 22.665 163.88 22.835 ;
      RECT 163.285 21.985 163.455 22.155 ;
      RECT 162.89 21.645 163.06 21.815 ;
      RECT 162.405 16.885 162.575 17.055 ;
      RECT 162.405 19.265 162.575 19.435 ;
      RECT 162.405 22.325 162.575 22.495 ;
      RECT 160.565 15.865 160.735 16.035 ;
      RECT 160.565 23.005 160.735 23.175 ;
      RECT 160.105 20.285 160.275 20.455 ;
      RECT 160.105 26.745 160.275 26.915 ;
      RECT 159.415 27.765 159.585 27.935 ;
      RECT 158.725 28.105 158.895 28.275 ;
      RECT 158.265 24.705 158.435 24.875 ;
      RECT 158.265 28.105 158.435 28.275 ;
      RECT 158.255 16.545 158.425 16.715 ;
      RECT 158.255 21.985 158.425 22.155 ;
      RECT 157.82 16.205 157.99 16.375 ;
      RECT 157.82 21.645 157.99 21.815 ;
      RECT 157.795 19.605 157.965 19.775 ;
      RECT 157.575 24.705 157.745 24.875 ;
      RECT 157.575 27.765 157.745 27.935 ;
      RECT 157.36 19.945 157.53 20.115 ;
      RECT 156.885 24.705 157.055 24.875 ;
      RECT 156.885 27.765 157.055 27.935 ;
      RECT 156.425 24.365 156.595 24.535 ;
      RECT 156.25 16.205 156.42 16.375 ;
      RECT 156.25 21.645 156.42 21.815 ;
      RECT 155.79 19.945 155.96 20.115 ;
      RECT 155.735 16.545 155.905 16.715 ;
      RECT 155.735 21.985 155.905 22.155 ;
      RECT 155.735 24.705 155.905 24.875 ;
      RECT 155.275 19.605 155.445 19.775 ;
      RECT 155.045 24.025 155.215 24.195 ;
      RECT 154.97 16.885 155.14 17.055 ;
      RECT 154.97 22.665 155.14 22.835 ;
      RECT 154.545 16.545 154.715 16.715 ;
      RECT 154.545 21.985 154.715 22.155 ;
      RECT 154.51 18.925 154.68 19.095 ;
      RECT 154.15 16.205 154.32 16.375 ;
      RECT 154.15 21.645 154.32 21.815 ;
      RECT 154.085 19.605 154.255 19.775 ;
      RECT 153.69 19.945 153.86 20.115 ;
      RECT 153.665 16.885 153.835 17.055 ;
      RECT 153.665 21.985 153.835 22.155 ;
      RECT 153.205 19.265 153.375 19.435 ;
      RECT 151.825 24.705 151.995 24.875 ;
      RECT 148.605 11.445 148.775 11.615 ;
      RECT 145.845 17.565 146.015 17.735 ;
      RECT 145.845 18.585 146.015 18.755 ;
      RECT 145.205 16.885 145.375 17.055 ;
      RECT 145.155 19.265 145.325 19.435 ;
      RECT 144.61 16.885 144.78 17.055 ;
      RECT 144.465 13.825 144.635 13.995 ;
      RECT 144.465 19.265 144.635 19.435 ;
      RECT 144.005 16.885 144.175 17.055 ;
      RECT 144.005 19.265 144.175 19.435 ;
      RECT 143.315 19.265 143.485 19.435 ;
      RECT 143.09 16.885 143.26 17.055 ;
      RECT 142.625 16.885 142.795 17.055 ;
      RECT 142.625 19.265 142.795 19.435 ;
      RECT 142.165 26.745 142.335 26.915 ;
      RECT 141.705 23.005 141.875 23.175 ;
      RECT 141.245 24.705 141.415 24.875 ;
      RECT 141.245 30.145 141.415 30.315 ;
      RECT 140.555 24.705 140.725 24.875 ;
      RECT 140.555 30.145 140.725 30.315 ;
      RECT 139.865 18.585 140.035 18.755 ;
      RECT 139.865 24.705 140.035 24.875 ;
      RECT 139.865 29.805 140.035 29.975 ;
      RECT 139.855 27.425 140.025 27.595 ;
      RECT 139.42 27.085 139.59 27.255 ;
      RECT 139.405 11.445 139.575 11.615 ;
      RECT 139.405 24.365 139.575 24.535 ;
      RECT 139.405 30.145 139.575 30.315 ;
      RECT 139.395 21.985 139.565 22.155 ;
      RECT 138.96 21.645 139.13 21.815 ;
      RECT 138.715 24.705 138.885 24.875 ;
      RECT 138.715 30.145 138.885 30.315 ;
      RECT 138.025 17.565 138.195 17.735 ;
      RECT 138.025 24.025 138.195 24.195 ;
      RECT 138.025 29.465 138.195 29.635 ;
      RECT 137.85 27.085 138.02 27.255 ;
      RECT 137.555 19.605 137.725 19.775 ;
      RECT 137.39 21.645 137.56 21.815 ;
      RECT 137.335 16.885 137.505 17.055 ;
      RECT 137.335 27.425 137.505 27.595 ;
      RECT 137.12 19.945 137.29 20.115 ;
      RECT 136.875 21.985 137.045 22.155 ;
      RECT 136.57 16.885 136.74 17.055 ;
      RECT 136.57 28.105 136.74 28.275 ;
      RECT 136.185 17.225 136.355 17.395 ;
      RECT 136.145 27.425 136.315 27.595 ;
      RECT 136.11 22.665 136.28 22.835 ;
      RECT 135.75 27.085 135.92 27.255 ;
      RECT 135.685 21.985 135.855 22.155 ;
      RECT 135.55 19.945 135.72 20.115 ;
      RECT 135.495 16.885 135.665 17.055 ;
      RECT 135.29 21.645 135.46 21.815 ;
      RECT 135.265 27.425 135.435 27.595 ;
      RECT 135.035 19.605 135.205 19.775 ;
      RECT 134.805 16.885 134.975 17.055 ;
      RECT 134.805 22.325 134.975 22.495 ;
      RECT 134.345 23.005 134.515 23.175 ;
      RECT 134.27 19.265 134.44 19.435 ;
      RECT 133.885 13.825 134.055 13.995 ;
      RECT 133.845 19.605 134.015 19.775 ;
      RECT 133.45 19.945 133.62 20.115 ;
      RECT 132.965 19.605 133.135 19.775 ;
      RECT 131.585 21.305 131.755 21.475 ;
      RECT 131.585 26.745 131.755 26.915 ;
      RECT 131.585 28.445 131.755 28.615 ;
      RECT 129.275 21.985 129.445 22.155 ;
      RECT 129.275 27.425 129.445 27.595 ;
      RECT 128.84 21.645 129.01 21.815 ;
      RECT 128.84 27.085 129.01 27.255 ;
      RECT 128.825 17.565 128.995 17.735 ;
      RECT 128.135 16.885 128.305 17.055 ;
      RECT 127.445 16.885 127.615 17.055 ;
      RECT 127.27 21.645 127.44 21.815 ;
      RECT 127.27 27.085 127.44 27.255 ;
      RECT 126.985 17.225 127.155 17.395 ;
      RECT 126.755 21.985 126.925 22.155 ;
      RECT 126.755 27.425 126.925 27.595 ;
      RECT 126.205 16.885 126.375 17.055 ;
      RECT 125.99 22.665 126.16 22.835 ;
      RECT 125.99 28.105 126.16 28.275 ;
      RECT 125.605 16.885 125.775 17.055 ;
      RECT 125.565 21.985 125.735 22.155 ;
      RECT 125.565 27.425 125.735 27.595 ;
      RECT 125.17 21.645 125.34 21.815 ;
      RECT 125.17 27.085 125.34 27.255 ;
      RECT 125.145 18.585 125.315 18.755 ;
      RECT 125.145 25.725 125.315 25.895 ;
      RECT 124.685 22.325 124.855 22.495 ;
      RECT 124.685 27.425 124.855 27.595 ;
      RECT 122.845 11.445 123.015 11.615 ;
      RECT 122.845 28.445 123.015 28.615 ;
      RECT 122.845 29.465 123.015 29.635 ;
      RECT 122.835 19.605 123.005 19.775 ;
      RECT 122.835 25.045 123.005 25.215 ;
      RECT 122.4 19.945 122.57 20.115 ;
      RECT 122.4 25.385 122.57 25.555 ;
      RECT 122.385 16.885 122.555 17.055 ;
      RECT 122.155 27.765 122.325 27.935 ;
      RECT 122.155 30.145 122.325 30.315 ;
      RECT 121.465 13.145 121.635 13.315 ;
      RECT 121.465 28.105 121.635 28.275 ;
      RECT 121.465 29.805 121.635 29.975 ;
      RECT 121.005 27.765 121.175 27.935 ;
      RECT 121.005 29.805 121.175 29.975 ;
      RECT 120.83 19.945 121 20.115 ;
      RECT 120.83 25.385 121 25.555 ;
      RECT 120.825 13.825 120.995 13.995 ;
      RECT 120.315 19.605 120.485 19.775 ;
      RECT 120.315 25.045 120.485 25.215 ;
      RECT 120.315 27.765 120.485 27.935 ;
      RECT 120.315 30.145 120.485 30.315 ;
      RECT 120.085 13.485 120.255 13.655 ;
      RECT 119.625 27.765 119.795 27.935 ;
      RECT 119.625 30.145 119.795 30.315 ;
      RECT 119.55 13.485 119.72 13.655 ;
      RECT 119.55 18.925 119.72 19.095 ;
      RECT 119.55 24.365 119.72 24.535 ;
      RECT 119.55 32.185 119.72 32.355 ;
      RECT 119.125 19.605 119.295 19.775 ;
      RECT 119.125 25.045 119.295 25.215 ;
      RECT 118.985 13.825 119.155 13.995 ;
      RECT 118.73 19.945 118.9 20.115 ;
      RECT 118.73 25.385 118.9 25.555 ;
      RECT 118.245 13.825 118.415 13.995 ;
      RECT 118.245 19.605 118.415 19.775 ;
      RECT 118.245 24.705 118.415 24.875 ;
      RECT 117.325 21.305 117.495 21.475 ;
      RECT 115.945 24.025 116.115 24.195 ;
      RECT 115.485 13.825 115.655 13.995 ;
      RECT 115.255 24.705 115.425 24.875 ;
      RECT 115.015 21.985 115.185 22.155 ;
      RECT 114.58 21.645 114.75 21.815 ;
      RECT 114.565 17.565 114.735 17.735 ;
      RECT 114.565 19.265 114.735 19.435 ;
      RECT 114.565 24.705 114.735 24.875 ;
      RECT 114.105 24.365 114.275 24.535 ;
      RECT 113.875 16.885 114.045 17.055 ;
      RECT 113.415 24.705 113.585 24.875 ;
      RECT 113.185 17.225 113.355 17.395 ;
      RECT 113.01 21.645 113.18 21.815 ;
      RECT 112.725 16.885 112.895 17.055 ;
      RECT 112.725 24.705 112.895 24.875 ;
      RECT 112.495 21.985 112.665 22.155 ;
      RECT 112.035 16.885 112.205 17.055 ;
      RECT 111.73 22.665 111.9 22.835 ;
      RECT 111.345 16.885 111.515 17.055 ;
      RECT 111.305 21.985 111.475 22.155 ;
      RECT 110.91 21.645 111.08 21.815 ;
      RECT 110.425 22.325 110.595 22.495 ;
      RECT 103.525 13.825 103.695 13.995 ;
      RECT 103.525 16.885 103.695 17.055 ;
      RECT 102.605 21.305 102.775 21.475 ;
      RECT 100.765 18.585 100.935 18.755 ;
      RECT 100.765 20.285 100.935 20.455 ;
      RECT 100.295 21.985 100.465 22.155 ;
      RECT 99.86 21.645 100.03 21.815 ;
      RECT 98.465 11.445 98.635 11.615 ;
      RECT 98.455 19.605 98.625 19.775 ;
      RECT 98.29 21.645 98.46 21.815 ;
      RECT 98.02 19.945 98.19 20.115 ;
      RECT 98.005 16.885 98.175 17.055 ;
      RECT 98.005 24.025 98.175 24.195 ;
      RECT 97.775 21.985 97.945 22.155 ;
      RECT 97.4 16.885 97.57 17.055 ;
      RECT 97.085 29.465 97.255 29.635 ;
      RECT 97.01 22.665 97.18 22.835 ;
      RECT 96.625 17.225 96.795 17.395 ;
      RECT 96.585 21.985 96.755 22.155 ;
      RECT 96.45 19.945 96.62 20.115 ;
      RECT 96.395 30.145 96.565 30.315 ;
      RECT 96.19 21.645 96.36 21.815 ;
      RECT 96.165 16.885 96.335 17.055 ;
      RECT 96.16 13.145 96.33 13.315 ;
      RECT 95.935 19.605 96.105 19.775 ;
      RECT 95.705 22.325 95.875 22.495 ;
      RECT 95.705 30.145 95.875 30.315 ;
      RECT 95.695 25.045 95.865 25.215 ;
      RECT 95.475 13.825 95.645 13.995 ;
      RECT 95.475 16.885 95.645 17.055 ;
      RECT 95.26 25.385 95.43 25.555 ;
      RECT 95.245 29.805 95.415 29.975 ;
      RECT 95.17 18.925 95.34 19.095 ;
      RECT 94.785 13.485 94.955 13.655 ;
      RECT 94.785 17.565 94.955 17.735 ;
      RECT 94.745 19.605 94.915 19.775 ;
      RECT 94.555 30.145 94.725 30.315 ;
      RECT 94.35 19.945 94.52 20.115 ;
      RECT 94.325 13.825 94.495 13.995 ;
      RECT 93.865 19.605 94.035 19.775 ;
      RECT 93.865 30.145 94.035 30.315 ;
      RECT 93.69 25.385 93.86 25.555 ;
      RECT 93.635 13.825 93.805 13.995 ;
      RECT 93.175 25.045 93.345 25.215 ;
      RECT 92.945 13.825 93.115 13.995 ;
      RECT 92.41 24.365 92.58 24.535 ;
      RECT 91.985 25.045 92.155 25.215 ;
      RECT 91.59 25.385 91.76 25.555 ;
      RECT 91.565 11.445 91.735 11.615 ;
      RECT 91.105 24.705 91.275 24.875 ;
      RECT 87.885 21.305 88.055 21.475 ;
      RECT 86.045 20.285 86.215 20.455 ;
      RECT 85.575 21.985 85.745 22.155 ;
      RECT 85.355 19.265 85.525 19.435 ;
      RECT 85.14 21.645 85.31 21.815 ;
      RECT 84.665 16.885 84.835 17.055 ;
      RECT 84.665 19.265 84.835 19.435 ;
      RECT 84.205 18.925 84.375 19.095 ;
      RECT 84.205 24.025 84.375 24.195 ;
      RECT 83.975 16.885 84.145 17.055 ;
      RECT 83.745 29.465 83.915 29.635 ;
      RECT 83.57 21.645 83.74 21.815 ;
      RECT 83.515 19.265 83.685 19.435 ;
      RECT 83.285 16.885 83.455 17.055 ;
      RECT 83.055 21.985 83.225 22.155 ;
      RECT 83.055 30.145 83.225 30.315 ;
      RECT 82.825 11.445 82.995 11.615 ;
      RECT 82.825 16.885 82.995 17.055 ;
      RECT 82.825 19.265 82.995 19.435 ;
      RECT 82.405 29.805 82.575 29.975 ;
      RECT 82.365 18.585 82.535 18.755 ;
      RECT 82.32 22.665 82.49 22.835 ;
      RECT 82.135 16.885 82.305 17.055 ;
      RECT 81.905 29.745 82.075 29.915 ;
      RECT 81.895 25.045 82.065 25.215 ;
      RECT 81.865 21.985 82.035 22.155 ;
      RECT 81.47 21.645 81.64 21.815 ;
      RECT 81.46 25.385 81.63 25.555 ;
      RECT 81.445 17.565 81.615 17.735 ;
      RECT 81.215 30.145 81.385 30.315 ;
      RECT 80.985 22.325 81.155 22.495 ;
      RECT 80.525 23.005 80.695 23.175 ;
      RECT 80.525 30.145 80.695 30.315 ;
      RECT 80.055 19.605 80.225 19.775 ;
      RECT 79.89 25.385 80.06 25.555 ;
      RECT 79.62 19.945 79.79 20.115 ;
      RECT 79.375 25.045 79.545 25.215 ;
      RECT 78.61 24.365 78.78 24.535 ;
      RECT 78.185 25.045 78.355 25.215 ;
      RECT 78.05 19.945 78.22 20.115 ;
      RECT 77.79 25.385 77.96 25.555 ;
      RECT 77.535 19.605 77.705 19.775 ;
      RECT 77.305 25.045 77.475 25.215 ;
      RECT 77.305 29.465 77.475 29.635 ;
      RECT 76.77 18.925 76.94 19.095 ;
      RECT 76.615 30.145 76.785 30.315 ;
      RECT 76.345 19.605 76.515 19.775 ;
      RECT 75.95 19.945 76.12 20.115 ;
      RECT 75.925 29.805 76.095 29.975 ;
      RECT 75.465 19.265 75.635 19.435 ;
      RECT 75.465 29.805 75.635 29.975 ;
      RECT 74.775 30.145 74.945 30.315 ;
      RECT 74.085 11.445 74.255 11.615 ;
      RECT 74.085 16.885 74.255 17.055 ;
      RECT 74.085 30.145 74.255 30.315 ;
      RECT 73.165 23.005 73.335 23.175 ;
      RECT 71.785 19.265 71.955 19.435 ;
      RECT 71.785 27.765 71.955 27.935 ;
      RECT 71.75 16.885 71.92 17.055 ;
      RECT 71.18 16.885 71.35 17.055 ;
      RECT 71.18 19.265 71.35 19.435 ;
      RECT 71.095 27.765 71.265 27.935 ;
      RECT 70.855 21.985 71.025 22.155 ;
      RECT 70.42 21.645 70.59 21.815 ;
      RECT 70.405 17.225 70.575 17.395 ;
      RECT 70.405 19.265 70.575 19.435 ;
      RECT 70.405 28.105 70.575 28.275 ;
      RECT 69.945 16.885 70.115 17.055 ;
      RECT 69.945 18.925 70.115 19.095 ;
      RECT 69.945 27.765 70.115 27.935 ;
      RECT 69.255 16.885 69.425 17.055 ;
      RECT 69.255 19.265 69.425 19.435 ;
      RECT 69.255 27.765 69.425 27.935 ;
      RECT 68.85 21.645 69.02 21.815 ;
      RECT 68.565 17.565 68.735 17.735 ;
      RECT 68.565 20.285 68.735 20.455 ;
      RECT 68.565 28.445 68.735 28.615 ;
      RECT 68.335 21.985 68.505 22.155 ;
      RECT 67.57 22.325 67.74 22.495 ;
      RECT 67.145 21.985 67.315 22.155 ;
      RECT 66.75 21.645 66.92 21.815 ;
      RECT 66.725 13.825 66.895 13.995 ;
      RECT 66.265 15.865 66.435 16.035 ;
      RECT 66.265 18.585 66.435 18.755 ;
      RECT 66.265 22.325 66.435 22.495 ;
      RECT 66.265 26.745 66.435 26.915 ;
      RECT 66.265 31.165 66.435 31.335 ;
      RECT 65.805 24.705 65.975 24.875 ;
      RECT 63.965 13.825 64.135 13.995 ;
      RECT 63.955 16.545 64.125 16.715 ;
      RECT 63.955 19.605 64.125 19.775 ;
      RECT 63.955 27.425 64.125 27.595 ;
      RECT 63.955 30.485 64.125 30.655 ;
      RECT 63.52 16.205 63.69 16.375 ;
      RECT 63.52 19.945 63.69 20.115 ;
      RECT 63.52 27.085 63.69 27.255 ;
      RECT 63.52 30.825 63.69 30.995 ;
      RECT 63.275 13.825 63.445 13.995 ;
      RECT 62.585 11.445 62.755 11.615 ;
      RECT 62.585 13.825 62.755 13.995 ;
      RECT 62.125 13.485 62.295 13.655 ;
      RECT 61.95 16.205 62.12 16.375 ;
      RECT 61.95 19.945 62.12 20.115 ;
      RECT 61.95 27.085 62.12 27.255 ;
      RECT 61.95 30.825 62.12 30.995 ;
      RECT 61.435 13.825 61.605 13.995 ;
      RECT 61.435 16.545 61.605 16.715 ;
      RECT 61.435 19.605 61.605 19.775 ;
      RECT 61.435 27.425 61.605 27.595 ;
      RECT 61.435 30.485 61.605 30.655 ;
      RECT 60.745 14.845 60.915 15.015 ;
      RECT 60.67 16.885 60.84 17.055 ;
      RECT 60.67 18.925 60.84 19.095 ;
      RECT 60.67 27.765 60.84 27.935 ;
      RECT 60.67 29.805 60.84 29.975 ;
      RECT 60.285 23.005 60.455 23.175 ;
      RECT 60.245 16.545 60.415 16.715 ;
      RECT 60.245 19.605 60.415 19.775 ;
      RECT 60.245 27.425 60.415 27.595 ;
      RECT 60.245 30.485 60.415 30.655 ;
      RECT 59.85 16.205 60.02 16.375 ;
      RECT 59.85 19.945 60.02 20.115 ;
      RECT 59.85 27.085 60.02 27.255 ;
      RECT 59.85 30.825 60.02 30.995 ;
      RECT 59.365 16.885 59.535 17.055 ;
      RECT 59.365 19.265 59.535 19.435 ;
      RECT 59.365 27.765 59.535 27.935 ;
      RECT 59.365 30.145 59.535 30.315 ;
      RECT 58.445 21.305 58.615 21.475 ;
      RECT 57.065 15.865 57.235 16.035 ;
      RECT 56.605 18.585 56.775 18.755 ;
      RECT 56.605 24.025 56.775 24.195 ;
      RECT 56.135 21.985 56.305 22.155 ;
      RECT 55.7 21.645 55.87 21.815 ;
      RECT 55.685 32.185 55.855 32.355 ;
      RECT 55.225 34.905 55.395 35.075 ;
      RECT 54.755 16.545 54.925 16.715 ;
      RECT 54.32 16.205 54.49 16.375 ;
      RECT 54.295 19.605 54.465 19.775 ;
      RECT 54.295 25.045 54.465 25.215 ;
      RECT 54.13 21.645 54.3 21.815 ;
      RECT 53.86 19.945 54.03 20.115 ;
      RECT 53.86 25.385 54.03 25.555 ;
      RECT 53.845 14.845 54.015 15.015 ;
      RECT 53.615 21.985 53.785 22.155 ;
      RECT 53.375 32.865 53.545 33.035 ;
      RECT 53.155 13.825 53.325 13.995 ;
      RECT 52.94 32.525 53.11 32.695 ;
      RECT 52.915 35.925 53.085 36.095 ;
      RECT 52.85 22.665 53.02 22.835 ;
      RECT 52.75 16.205 52.92 16.375 ;
      RECT 52.48 36.265 52.65 36.435 ;
      RECT 52.465 13.485 52.635 13.655 ;
      RECT 52.425 21.985 52.595 22.155 ;
      RECT 52.29 19.945 52.46 20.115 ;
      RECT 52.29 25.385 52.46 25.555 ;
      RECT 52.235 16.545 52.405 16.715 ;
      RECT 52.03 21.645 52.2 21.815 ;
      RECT 52.005 13.485 52.175 13.655 ;
      RECT 51.775 19.605 51.945 19.775 ;
      RECT 51.775 25.045 51.945 25.215 ;
      RECT 51.545 22.325 51.715 22.495 ;
      RECT 51.47 16.885 51.64 17.055 ;
      RECT 51.37 32.525 51.54 32.695 ;
      RECT 51.09 13.825 51.26 13.995 ;
      RECT 51.045 16.545 51.215 16.715 ;
      RECT 51.01 18.925 51.18 19.095 ;
      RECT 51.01 24.365 51.18 24.535 ;
      RECT 50.91 36.265 51.08 36.435 ;
      RECT 50.855 32.865 51.025 33.035 ;
      RECT 50.655 13.825 50.825 13.995 ;
      RECT 50.65 16.205 50.82 16.375 ;
      RECT 50.585 19.605 50.755 19.775 ;
      RECT 50.585 25.045 50.755 25.215 ;
      RECT 50.395 35.925 50.565 36.095 ;
      RECT 50.19 19.945 50.36 20.115 ;
      RECT 50.19 25.385 50.36 25.555 ;
      RECT 50.165 16.885 50.335 17.055 ;
      RECT 50.09 33.205 50.26 33.375 ;
      RECT 49.705 19.265 49.875 19.435 ;
      RECT 49.705 24.705 49.875 24.875 ;
      RECT 49.665 32.865 49.835 33.035 ;
      RECT 49.63 35.245 49.8 35.415 ;
      RECT 49.27 32.525 49.44 32.695 ;
      RECT 49.245 23.005 49.415 23.175 ;
      RECT 49.245 28.445 49.415 28.615 ;
      RECT 49.245 31.165 49.415 31.335 ;
      RECT 49.205 35.925 49.375 36.095 ;
      RECT 48.81 36.265 48.98 36.435 ;
      RECT 48.785 11.445 48.955 11.615 ;
      RECT 48.785 32.865 48.955 33.035 ;
      RECT 48.555 22.325 48.725 22.495 ;
      RECT 48.555 27.765 48.725 27.935 ;
      RECT 48.555 30.145 48.725 30.315 ;
      RECT 48.325 35.925 48.495 36.095 ;
      RECT 47.865 17.565 48.035 17.735 ;
      RECT 47.865 22.325 48.035 22.495 ;
      RECT 47.865 28.105 48.035 28.275 ;
      RECT 47.865 29.805 48.035 29.975 ;
      RECT 47.405 14.845 47.575 15.015 ;
      RECT 47.405 22.665 47.575 22.835 ;
      RECT 47.405 30.145 47.575 30.315 ;
      RECT 47.175 16.885 47.345 17.055 ;
      RECT 47.175 27.765 47.345 27.935 ;
      RECT 46.715 22.325 46.885 22.495 ;
      RECT 46.715 27.765 46.885 27.935 ;
      RECT 46.715 30.145 46.885 30.315 ;
      RECT 46.485 16.885 46.655 17.055 ;
      RECT 46.025 13.825 46.195 13.995 ;
      RECT 46.025 17.225 46.195 17.395 ;
      RECT 46.025 22.325 46.195 22.495 ;
      RECT 46.025 27.765 46.195 27.935 ;
      RECT 46.025 30.145 46.195 30.315 ;
      RECT 45.59 13.825 45.76 13.995 ;
      RECT 45.565 14.845 45.735 15.015 ;
      RECT 45.335 16.885 45.505 17.055 ;
      RECT 44.645 16.885 44.815 17.055 ;
      RECT 40.505 16.885 40.675 17.055 ;
      RECT 40.505 27.765 40.675 27.935 ;
      RECT 37.745 13.825 37.915 13.995 ;
      RECT 30.845 11.445 31.015 11.615 ;
      RECT 30.845 16.885 31.015 17.055 ;
      RECT 22.105 24.705 22.275 24.875 ;
      RECT 20.265 13.825 20.435 13.995 ;
      RECT 20.265 16.885 20.435 17.055 ;
    LAYER met1 ;
      RECT 176.68 13.84 183.26 13.98 ;
      RECT 183.12 13.5 183.26 13.98 ;
      RECT 176.68 13.5 176.82 13.98 ;
      RECT 183.95 13.44 184.27 13.7 ;
      RECT 167.39 13.44 167.71 13.7 ;
      RECT 169.245 13.455 169.535 13.685 ;
      RECT 183.12 13.5 184.27 13.64 ;
      RECT 173.46 13.5 176.82 13.64 ;
      RECT 167.39 13.5 170.38 13.64 ;
      RECT 170.24 13.33 170.38 13.64 ;
      RECT 173.46 13.33 173.6 13.64 ;
      RECT 170.24 13.33 173.6 13.47 ;
      RECT 181.655 21.955 181.945 22.185 ;
      RECT 179.135 21.955 179.425 22.185 ;
      RECT 177.945 21.955 178.235 22.185 ;
      RECT 177.945 22 181.945 22.14 ;
      RECT 181.22 21.615 181.51 21.845 ;
      RECT 179.65 21.615 179.94 21.845 ;
      RECT 177.55 21.615 177.84 21.845 ;
      RECT 177.55 21.66 181.51 21.8 ;
      RECT 131.525 28.415 131.815 28.645 ;
      RECT 155.52 28.46 158.88 28.6 ;
      RECT 158.74 28.075 158.88 28.6 ;
      RECT 135.74 28.46 138.18 28.6 ;
      RECT 138.04 28.12 138.18 28.6 ;
      RECT 131.525 28.46 132.66 28.6 ;
      RECT 132.52 28.29 132.66 28.6 ;
      RECT 155.52 28.29 155.66 28.6 ;
      RECT 135.74 28.29 135.88 28.6 ;
      RECT 150 28.29 155.66 28.43 ;
      RECT 132.52 28.29 135.88 28.43 ;
      RECT 181.19 28.06 181.51 28.32 ;
      RECT 158.665 28.075 158.955 28.305 ;
      RECT 150 28.12 150.14 28.43 ;
      RECT 180.36 28.12 181.51 28.26 ;
      RECT 158.665 28.12 168.54 28.26 ;
      RECT 168.4 27.78 168.54 28.26 ;
      RECT 138.04 28.12 150.14 28.26 ;
      RECT 180.36 27.78 180.5 28.26 ;
      RECT 168.4 27.78 180.5 27.92 ;
      RECT 175.67 22.62 175.99 22.88 ;
      RECT 178.37 22.635 178.66 22.865 ;
      RECT 175.67 22.68 178.66 22.82 ;
      RECT 175.67 16.84 175.99 17.1 ;
      RECT 177.065 16.855 177.355 17.085 ;
      RECT 175.67 16.9 177.355 17.04 ;
      RECT 177.065 21.955 177.355 22.185 ;
      RECT 172.54 22 177.355 22.14 ;
      RECT 172.54 21.66 172.68 22.14 ;
      RECT 170.15 21.6 170.47 21.86 ;
      RECT 171.085 21.615 171.375 21.845 ;
      RECT 170.15 21.66 172.68 21.8 ;
      RECT 175.67 15.82 175.99 16.08 ;
      RECT 176.145 15.835 176.435 16.065 ;
      RECT 175.67 15.88 176.435 16.02 ;
      RECT 175.67 14.46 175.99 14.72 ;
      RECT 158.28 14.52 175.99 14.66 ;
      RECT 169.78 13.795 169.92 14.66 ;
      RECT 158.28 14.18 158.42 14.66 ;
      RECT 148.62 14.18 158.42 14.32 ;
      RECT 148.62 13.84 148.76 14.32 ;
      RECT 145.31 13.78 145.63 14.04 ;
      RECT 169.705 13.795 169.995 14.025 ;
      RECT 144.405 13.795 144.695 14.025 ;
      RECT 144.405 13.84 148.76 13.98 ;
      RECT 175.67 21.26 175.99 21.52 ;
      RECT 169.245 21.275 169.535 21.505 ;
      RECT 169.245 21.32 175.99 21.46 ;
      RECT 169.245 24.335 169.535 24.565 ;
      RECT 169.245 24.38 175.9 24.52 ;
      RECT 175.76 23.98 175.9 24.52 ;
      RECT 175.67 23.98 175.99 24.24 ;
      RECT 167.39 20.24 167.71 20.5 ;
      RECT 173.845 20.255 174.135 20.485 ;
      RECT 167.39 20.3 174.135 20.44 ;
      RECT 173.835 16.515 174.125 16.745 ;
      RECT 171.315 16.515 171.605 16.745 ;
      RECT 170.125 16.515 170.415 16.745 ;
      RECT 170.125 16.56 174.125 16.7 ;
      RECT 173.4 16.175 173.69 16.405 ;
      RECT 171.83 16.175 172.12 16.405 ;
      RECT 169.73 16.175 170.02 16.405 ;
      RECT 169.73 16.22 173.69 16.36 ;
      RECT 148.07 11.4 148.39 11.66 ;
      RECT 148.545 11.415 148.835 11.645 ;
      RECT 148.07 11.46 148.835 11.6 ;
      RECT 148.62 10.44 148.76 11.645 ;
      RECT 166.1 11.12 172.22 11.26 ;
      RECT 172.08 10.44 172.22 11.26 ;
      RECT 154.6 11.12 161.18 11.26 ;
      RECT 161.04 10.61 161.18 11.26 ;
      RECT 166.1 10.61 166.24 11.26 ;
      RECT 154.6 10.61 154.74 11.26 ;
      RECT 161.04 10.61 166.24 10.75 ;
      RECT 149.54 10.61 154.74 10.75 ;
      RECT 172.91 10.38 173.23 10.64 ;
      RECT 149.54 10.44 149.68 10.75 ;
      RECT 172.08 10.44 173.23 10.58 ;
      RECT 148.62 10.44 149.68 10.58 ;
      RECT 172.91 19.9 173.23 20.16 ;
      RECT 172.465 19.915 172.755 20.145 ;
      RECT 172.465 19.96 173.23 20.1 ;
      RECT 172.91 23.98 173.23 24.24 ;
      RECT 171.085 23.995 171.375 24.225 ;
      RECT 171.085 24.04 173.23 24.18 ;
      RECT 167.39 25.34 167.71 25.6 ;
      RECT 167.39 25.4 171.76 25.54 ;
      RECT 171.62 24.675 171.76 25.54 ;
      RECT 172.91 24.66 173.23 24.92 ;
      RECT 171.545 24.675 171.835 24.905 ;
      RECT 171.545 24.72 173.23 24.86 ;
      RECT 145.31 17.52 145.63 17.78 ;
      RECT 168.86 17.58 171.3 17.72 ;
      RECT 171.16 16.9 171.3 17.72 ;
      RECT 168.86 17.24 169 17.72 ;
      RECT 153.22 17.41 163.02 17.55 ;
      RECT 162.88 17.24 163.02 17.55 ;
      RECT 145.4 17.24 145.54 17.78 ;
      RECT 153.22 17.24 153.36 17.55 ;
      RECT 162.88 17.24 169 17.38 ;
      RECT 145.4 17.24 153.36 17.38 ;
      RECT 170.58 16.855 170.87 17.085 ;
      RECT 170.58 16.9 171.3 17.04 ;
      RECT 170.15 17.18 170.47 17.44 ;
      RECT 170.24 16.9 170.38 17.44 ;
      RECT 169.245 16.855 169.535 17.085 ;
      RECT 169.245 16.9 170.38 17.04 ;
      RECT 150.83 25.68 151.15 25.94 ;
      RECT 150 25.74 158.42 25.88 ;
      RECT 158.28 24.675 158.42 25.88 ;
      RECT 150 25.4 150.14 25.88 ;
      RECT 143.1 25.4 150.14 25.54 ;
      RECT 143.1 24.72 143.24 25.54 ;
      RECT 159.2 25.06 165.32 25.2 ;
      RECT 165.18 24.72 165.32 25.2 ;
      RECT 159.2 24.72 159.34 25.2 ;
      RECT 142.55 24.66 142.87 24.92 ;
      RECT 170.165 24.675 170.455 24.905 ;
      RECT 158.205 24.675 158.495 24.905 ;
      RECT 141.185 24.675 141.475 24.905 ;
      RECT 165.18 24.72 170.455 24.86 ;
      RECT 158.205 24.72 159.34 24.86 ;
      RECT 141.185 24.72 143.24 24.86 ;
      RECT 167.48 24.32 167.62 24.86 ;
      RECT 167.39 24.32 167.71 24.58 ;
      RECT 170.155 19.575 170.445 19.805 ;
      RECT 167.635 19.575 167.925 19.805 ;
      RECT 166.445 19.575 166.735 19.805 ;
      RECT 166.445 19.62 170.445 19.76 ;
      RECT 169.72 19.915 170.01 20.145 ;
      RECT 168.15 19.915 168.44 20.145 ;
      RECT 166.05 19.915 166.34 20.145 ;
      RECT 166.05 19.96 170.01 20.1 ;
      RECT 164.63 22.96 164.95 23.22 ;
      RECT 169.245 22.975 169.535 23.205 ;
      RECT 168.4 23.02 169.535 23.16 ;
      RECT 164.63 23.02 165.78 23.16 ;
      RECT 165.64 22.68 165.78 23.16 ;
      RECT 168.4 22.68 168.54 23.16 ;
      RECT 165.64 22.68 168.54 22.82 ;
      RECT 159.11 13.78 159.43 14.04 ;
      RECT 168.555 13.795 168.845 14.025 ;
      RECT 159.11 13.84 168.845 13.98 ;
      RECT 167.39 14.8 167.71 15.06 ;
      RECT 167.865 14.815 168.155 15.045 ;
      RECT 167.39 14.86 168.155 15 ;
      RECT 167.39 12.08 167.71 12.34 ;
      RECT 164.26 12.14 167.71 12.28 ;
      RECT 164.26 11.415 164.4 12.28 ;
      RECT 164.185 11.415 164.475 11.645 ;
      RECT 162.345 19.235 162.635 19.465 ;
      RECT 162.345 19.28 164.4 19.42 ;
      RECT 164.26 18.6 164.4 19.42 ;
      RECT 167.39 18.54 167.71 18.8 ;
      RECT 164.26 18.6 167.71 18.74 ;
      RECT 157.515 27.735 157.805 27.965 ;
      RECT 157.59 27.1 157.73 27.965 ;
      RECT 143.56 27.44 150.14 27.58 ;
      RECT 150 27.1 150.14 27.58 ;
      RECT 143.56 27.1 143.7 27.58 ;
      RECT 142.55 27.04 142.87 27.3 ;
      RECT 150 27.1 167.62 27.24 ;
      RECT 167.48 26.7 167.62 27.24 ;
      RECT 142.55 27.1 143.7 27.24 ;
      RECT 153.68 26.7 153.82 27.24 ;
      RECT 167.39 26.7 167.71 26.96 ;
      RECT 153.59 26.7 153.91 26.96 ;
      RECT 166.935 21.955 167.225 22.185 ;
      RECT 164.415 21.955 164.705 22.185 ;
      RECT 163.225 21.955 163.515 22.185 ;
      RECT 163.225 22 167.225 22.14 ;
      RECT 166.87 18.895 167.16 19.125 ;
      RECT 165.105 18.895 165.395 19.125 ;
      RECT 165.105 18.94 167.16 19.08 ;
      RECT 166.5 21.615 166.79 21.845 ;
      RECT 164.93 21.615 165.22 21.845 ;
      RECT 162.83 21.615 163.12 21.845 ;
      RECT 162.83 21.66 166.79 21.8 ;
      RECT 164.63 19.22 164.95 19.48 ;
      RECT 165.565 19.235 165.855 19.465 ;
      RECT 164.63 19.28 165.855 19.42 ;
      RECT 156.365 24.335 156.655 24.565 ;
      RECT 160.12 24.38 163.94 24.52 ;
      RECT 163.8 24.04 163.94 24.52 ;
      RECT 160.12 24.21 160.26 24.52 ;
      RECT 157.36 24.21 160.26 24.35 ;
      RECT 156.44 24.04 156.58 24.565 ;
      RECT 164.63 23.98 164.95 24.24 ;
      RECT 157.36 24.04 157.5 24.35 ;
      RECT 163.8 24.04 164.95 24.18 ;
      RECT 156.44 24.04 157.5 24.18 ;
      RECT 161.87 22.96 162.19 23.22 ;
      RECT 161.96 22.68 162.1 23.22 ;
      RECT 163.65 22.635 163.94 22.865 ;
      RECT 161.96 22.68 163.94 22.82 ;
      RECT 156.35 16.84 156.67 17.1 ;
      RECT 162.345 16.855 162.635 17.085 ;
      RECT 161.5 16.9 162.635 17.04 ;
      RECT 156.35 16.9 159.34 17.04 ;
      RECT 159.2 16.56 159.34 17.04 ;
      RECT 161.5 16.56 161.64 17.04 ;
      RECT 159.2 16.56 161.64 16.7 ;
      RECT 161.87 22.28 162.19 22.54 ;
      RECT 162.345 22.295 162.635 22.525 ;
      RECT 161.87 22.34 162.635 22.48 ;
      RECT 161.87 26.7 162.19 26.96 ;
      RECT 160.045 26.715 160.335 26.945 ;
      RECT 160.045 26.76 162.19 26.9 ;
      RECT 143.945 16.855 144.235 17.085 ;
      RECT 127.385 16.855 127.675 17.085 ;
      RECT 144.02 15.88 144.16 17.085 ;
      RECT 127.46 15.88 127.6 17.085 ;
      RECT 125.99 16.16 126.31 16.42 ;
      RECT 146.32 16.22 150.14 16.36 ;
      RECT 150 16.05 150.14 16.36 ;
      RECT 137.12 16.22 141.86 16.36 ;
      RECT 141.72 15.88 141.86 16.36 ;
      RECT 125.99 16.22 127.6 16.36 ;
      RECT 146.32 15.88 146.46 16.36 ;
      RECT 137.12 16.05 137.26 16.36 ;
      RECT 150 16.05 153.36 16.19 ;
      RECT 153.22 15.88 153.36 16.19 ;
      RECT 133.44 16.05 137.26 16.19 ;
      RECT 160.505 15.835 160.795 16.065 ;
      RECT 133.44 15.88 133.58 16.19 ;
      RECT 153.22 15.88 160.795 16.02 ;
      RECT 141.72 15.88 146.46 16.02 ;
      RECT 127.46 15.88 133.58 16.02 ;
      RECT 156.35 22.96 156.67 23.22 ;
      RECT 160.505 22.975 160.795 23.205 ;
      RECT 156.35 23.02 160.795 23.16 ;
      RECT 134.27 20.24 134.59 20.5 ;
      RECT 160.045 20.255 160.335 20.485 ;
      RECT 152.3 20.3 160.335 20.44 ;
      RECT 141.72 20.3 145.08 20.44 ;
      RECT 144.94 20.13 145.08 20.44 ;
      RECT 134.27 20.3 138.64 20.44 ;
      RECT 138.5 19.96 138.64 20.44 ;
      RECT 152.3 19.96 152.44 20.44 ;
      RECT 144.02 19.235 144.16 20.44 ;
      RECT 141.72 19.96 141.86 20.44 ;
      RECT 144.94 20.13 149.22 20.27 ;
      RECT 149.08 19.96 149.22 20.27 ;
      RECT 149.08 19.96 152.44 20.1 ;
      RECT 138.5 19.96 141.86 20.1 ;
      RECT 143.945 19.235 144.235 19.465 ;
      RECT 159.11 27.72 159.43 27.98 ;
      RECT 159.11 27.735 159.645 27.965 ;
      RECT 159.11 22.28 159.43 22.54 ;
      RECT 148.07 22.28 148.39 22.54 ;
      RECT 148.07 22.34 159.43 22.48 ;
      RECT 156.35 28.06 156.67 28.32 ;
      RECT 158.205 28.075 158.495 28.305 ;
      RECT 156.35 28.12 158.495 28.26 ;
      RECT 158.195 16.515 158.485 16.745 ;
      RECT 155.675 16.515 155.965 16.745 ;
      RECT 154.485 16.515 154.775 16.745 ;
      RECT 154.485 16.56 158.485 16.7 ;
      RECT 158.195 21.955 158.485 22.185 ;
      RECT 155.675 21.955 155.965 22.185 ;
      RECT 154.485 21.955 154.775 22.185 ;
      RECT 154.485 22 158.485 22.14 ;
      RECT 157.76 16.175 158.05 16.405 ;
      RECT 156.19 16.175 156.48 16.405 ;
      RECT 154.09 16.175 154.38 16.405 ;
      RECT 154.09 16.22 158.05 16.36 ;
      RECT 157.76 21.615 158.05 21.845 ;
      RECT 156.19 21.615 156.48 21.845 ;
      RECT 154.09 21.615 154.38 21.845 ;
      RECT 154.09 21.66 158.05 21.8 ;
      RECT 157.735 19.575 158.025 19.805 ;
      RECT 155.215 19.575 155.505 19.805 ;
      RECT 154.025 19.575 154.315 19.805 ;
      RECT 154.025 19.62 158.025 19.76 ;
      RECT 153.59 25.34 153.91 25.6 ;
      RECT 153.59 25.4 157.04 25.54 ;
      RECT 156.9 25.06 157.04 25.54 ;
      RECT 156.9 25.06 157.73 25.2 ;
      RECT 157.59 24.675 157.73 25.2 ;
      RECT 157.515 24.675 157.805 24.905 ;
      RECT 157.3 19.915 157.59 20.145 ;
      RECT 155.73 19.915 156.02 20.145 ;
      RECT 153.63 19.915 153.92 20.145 ;
      RECT 153.63 19.96 157.59 20.1 ;
      RECT 154.6 25.06 156.58 25.2 ;
      RECT 156.44 24.72 156.58 25.2 ;
      RECT 154.6 24.72 154.74 25.2 ;
      RECT 156.825 24.675 157.115 24.905 ;
      RECT 151.765 24.675 152.055 24.905 ;
      RECT 156.44 24.72 157.115 24.86 ;
      RECT 148.62 24.72 154.74 24.86 ;
      RECT 148.62 24.38 148.76 24.86 ;
      RECT 145.31 24.32 145.63 24.58 ;
      RECT 139.345 24.335 139.635 24.565 ;
      RECT 139.345 24.38 148.76 24.52 ;
      RECT 150.83 27.72 151.15 27.98 ;
      RECT 156.825 27.735 157.115 27.965 ;
      RECT 150.83 27.78 157.115 27.92 ;
      RECT 140.8 30.67 143.7 30.81 ;
      RECT 143.56 30.5 143.7 30.81 ;
      RECT 140.8 30.5 140.94 30.81 ;
      RECT 143.56 30.5 156.58 30.64 ;
      RECT 156.44 30.1 156.58 30.64 ;
      RECT 139.88 30.5 140.94 30.64 ;
      RECT 139.88 30.16 140.02 30.64 ;
      RECT 156.35 30.1 156.67 30.36 ;
      RECT 139.345 30.115 139.635 30.345 ;
      RECT 139.345 30.16 140.02 30.3 ;
      RECT 137.03 24.66 137.35 24.92 ;
      RECT 155.675 24.675 155.965 24.905 ;
      RECT 138.655 24.675 138.945 24.905 ;
      RECT 136.66 24.72 138.945 24.86 ;
      RECT 138.04 24.38 138.18 24.86 ;
      RECT 136.66 24.38 136.8 24.86 ;
      RECT 155.75 24.38 155.89 24.905 ;
      RECT 152.3 24.38 155.89 24.52 ;
      RECT 138.04 24.38 139.1 24.52 ;
      RECT 138.96 24.04 139.1 24.52 ;
      RECT 128.84 24.38 136.8 24.52 ;
      RECT 152.3 24.21 152.44 24.52 ;
      RECT 128.84 23.98 128.98 24.52 ;
      RECT 149.54 24.21 152.44 24.35 ;
      RECT 148.07 23.98 148.39 24.24 ;
      RECT 128.75 23.98 129.07 24.24 ;
      RECT 149.54 24.04 149.68 24.35 ;
      RECT 138.96 24.04 149.68 24.18 ;
      RECT 153.59 23.98 153.91 24.24 ;
      RECT 154.985 23.995 155.275 24.225 ;
      RECT 153.59 24.04 155.275 24.18 ;
      RECT 154.91 16.855 155.2 17.085 ;
      RECT 154.14 16.9 155.2 17.04 ;
      RECT 154.14 16.56 154.28 17.04 ;
      RECT 150.83 16.5 151.15 16.76 ;
      RECT 150.83 16.56 154.28 16.7 ;
      RECT 153.59 22.62 153.91 22.88 ;
      RECT 154.91 22.635 155.2 22.865 ;
      RECT 153.59 22.68 155.2 22.82 ;
      RECT 149.08 19.28 152.44 19.42 ;
      RECT 152.3 18.94 152.44 19.42 ;
      RECT 149.08 18.94 149.22 19.42 ;
      RECT 148.07 18.88 148.39 19.14 ;
      RECT 154.45 18.895 154.74 19.125 ;
      RECT 152.3 18.94 154.74 19.08 ;
      RECT 148.07 18.94 149.22 19.08 ;
      RECT 153.59 19.22 153.91 19.48 ;
      RECT 153.145 19.235 153.435 19.465 ;
      RECT 153.145 19.28 153.91 19.42 ;
      RECT 141.185 30.115 141.475 30.345 ;
      RECT 141.185 30.16 143.24 30.3 ;
      RECT 143.1 29.82 143.24 30.3 ;
      RECT 150.83 29.76 151.15 30.02 ;
      RECT 143.1 29.82 151.15 29.96 ;
      RECT 148.07 16.84 148.39 17.1 ;
      RECT 145.145 16.855 145.435 17.085 ;
      RECT 145.145 16.9 148.39 17.04 ;
      RECT 148.07 17.52 148.39 17.78 ;
      RECT 145.785 17.535 146.075 17.765 ;
      RECT 145.785 17.58 148.39 17.72 ;
      RECT 148.07 19.56 148.39 19.82 ;
      RECT 144.48 19.62 148.39 19.76 ;
      RECT 144.48 19.235 144.62 19.76 ;
      RECT 144.405 19.235 144.695 19.465 ;
      RECT 145.31 18.54 145.63 18.8 ;
      RECT 145.785 18.555 146.075 18.785 ;
      RECT 145.31 18.6 146.075 18.74 ;
      RECT 144.55 16.855 144.84 17.085 ;
      RECT 144.625 16.22 144.765 17.085 ;
      RECT 145.31 16.16 145.63 16.42 ;
      RECT 144.625 16.22 145.63 16.36 ;
      RECT 145.31 26.7 145.63 26.96 ;
      RECT 142.105 26.715 142.395 26.945 ;
      RECT 142.105 26.76 145.63 26.9 ;
      RECT 145.095 19.235 145.385 19.465 ;
      RECT 145.17 18.94 145.31 19.465 ;
      RECT 142.64 18.94 145.31 19.08 ;
      RECT 142.64 18.54 142.78 19.08 ;
      RECT 142.55 18.54 142.87 18.8 ;
      RECT 142.55 19.9 142.87 20.16 ;
      RECT 142.64 19.62 142.78 20.16 ;
      RECT 142.64 19.62 143.47 19.76 ;
      RECT 143.33 19.235 143.47 19.76 ;
      RECT 143.255 19.235 143.545 19.465 ;
      RECT 143.03 16.855 143.32 17.085 ;
      RECT 143.105 16.56 143.245 17.085 ;
      RECT 142.64 16.56 143.245 16.7 ;
      RECT 142.64 16.16 142.78 16.7 ;
      RECT 142.55 16.16 142.87 16.42 ;
      RECT 142.55 17.52 142.87 17.78 ;
      RECT 142.18 17.58 142.87 17.72 ;
      RECT 142.18 16.9 142.32 17.72 ;
      RECT 137.275 16.855 137.565 17.085 ;
      RECT 137.275 16.9 142.32 17.04 ;
      RECT 142.55 19.22 142.87 19.48 ;
      RECT 138.04 19.28 142.87 19.42 ;
      RECT 138.04 19.11 138.18 19.42 ;
      RECT 135.28 19.11 138.18 19.25 ;
      RECT 135.28 18.6 135.42 19.25 ;
      RECT 128.75 18.54 129.07 18.8 ;
      RECT 128.75 18.6 135.42 18.74 ;
      RECT 142.55 25.34 142.87 25.6 ;
      RECT 140.57 25.4 142.87 25.54 ;
      RECT 140.57 24.675 140.71 25.54 ;
      RECT 140.495 24.675 140.785 24.905 ;
      RECT 140.495 30.115 140.785 30.345 ;
      RECT 140.57 29.48 140.71 30.345 ;
      RECT 142.55 29.42 142.87 29.68 ;
      RECT 140.57 29.48 142.87 29.62 ;
      RECT 142.55 31.12 142.87 31.38 ;
      RECT 139.88 31.18 142.87 31.32 ;
      RECT 139.88 31.01 140.02 31.32 ;
      RECT 137.12 31.01 140.02 31.15 ;
      RECT 137.12 30.5 137.26 31.15 ;
      RECT 121.48 30.84 123.92 30.98 ;
      RECT 123.78 30.5 123.92 30.98 ;
      RECT 121.48 30.16 121.62 30.98 ;
      RECT 125.99 30.44 126.31 30.7 ;
      RECT 123.78 30.5 137.26 30.64 ;
      RECT 120.47 30.1 120.79 30.36 ;
      RECT 120.255 30.115 120.79 30.345 ;
      RECT 120.255 30.16 121.62 30.3 ;
      RECT 139.79 22.96 140.11 23.22 ;
      RECT 141.645 22.975 141.935 23.205 ;
      RECT 139.79 23.02 141.935 23.16 ;
      RECT 139.79 11.4 140.11 11.66 ;
      RECT 139.345 11.415 139.635 11.645 ;
      RECT 139.345 11.46 140.11 11.6 ;
      RECT 139.79 17.52 140.11 17.78 ;
      RECT 137.965 17.535 138.255 17.765 ;
      RECT 137.965 17.58 140.11 17.72 ;
      RECT 124.24 29.99 126.68 30.13 ;
      RECT 126.54 29.82 126.68 30.13 ;
      RECT 139.79 29.76 140.11 30.02 ;
      RECT 121.405 29.775 121.695 30.005 ;
      RECT 124.24 29.82 124.38 30.13 ;
      RECT 126.54 29.82 138.64 29.96 ;
      RECT 138.5 29.48 138.64 29.96 ;
      RECT 121.405 29.82 124.38 29.96 ;
      RECT 139.88 29.48 140.02 30.02 ;
      RECT 138.5 29.48 140.02 29.62 ;
      RECT 137.03 18.54 137.35 18.8 ;
      RECT 139.805 18.555 140.095 18.785 ;
      RECT 137.03 18.6 140.095 18.74 ;
      RECT 136.2 25.4 139.1 25.54 ;
      RECT 138.96 25.06 139.1 25.54 ;
      RECT 136.2 25.06 136.34 25.54 ;
      RECT 131.51 25 131.83 25.26 ;
      RECT 138.96 25.06 140.02 25.2 ;
      RECT 139.88 24.675 140.02 25.2 ;
      RECT 131.51 25.06 136.34 25.2 ;
      RECT 139.805 24.675 140.095 24.905 ;
      RECT 139.795 27.395 140.085 27.625 ;
      RECT 137.275 27.395 137.565 27.625 ;
      RECT 136.085 27.395 136.375 27.625 ;
      RECT 136.085 27.44 140.085 27.58 ;
      RECT 139.36 27.055 139.65 27.285 ;
      RECT 137.79 27.055 138.08 27.285 ;
      RECT 135.69 27.055 135.98 27.285 ;
      RECT 135.69 27.1 139.65 27.24 ;
      RECT 139.335 21.955 139.625 22.185 ;
      RECT 136.815 21.955 137.105 22.185 ;
      RECT 135.625 21.955 135.915 22.185 ;
      RECT 135.625 22 139.625 22.14 ;
      RECT 138.9 21.615 139.19 21.845 ;
      RECT 137.33 21.615 137.62 21.845 ;
      RECT 135.23 21.615 135.52 21.845 ;
      RECT 135.23 21.66 139.19 21.8 ;
      RECT 137.03 30.1 137.35 30.36 ;
      RECT 138.655 30.115 138.945 30.345 ;
      RECT 137.03 30.16 138.945 30.3 ;
      RECT 137.03 23.98 137.35 24.24 ;
      RECT 137.965 23.995 138.255 24.225 ;
      RECT 137.03 24.04 138.255 24.18 ;
      RECT 137.03 29.42 137.35 29.68 ;
      RECT 137.965 29.435 138.255 29.665 ;
      RECT 137.03 29.48 138.255 29.62 ;
      RECT 137.495 19.575 137.785 19.805 ;
      RECT 134.975 19.575 135.265 19.805 ;
      RECT 133.785 19.575 134.075 19.805 ;
      RECT 133.785 19.62 137.785 19.76 ;
      RECT 137.03 13.44 137.35 13.7 ;
      RECT 123.23 13.44 123.55 13.7 ;
      RECT 120.025 13.455 120.315 13.685 ;
      RECT 129.3 13.5 137.35 13.64 ;
      RECT 120.025 13.5 124.38 13.64 ;
      RECT 124.24 13.33 124.38 13.64 ;
      RECT 129.3 13.33 129.44 13.64 ;
      RECT 124.24 13.33 129.44 13.47 ;
      RECT 137.03 17.52 137.35 17.78 ;
      RECT 136.2 17.58 137.35 17.72 ;
      RECT 136.2 17.195 136.34 17.72 ;
      RECT 136.125 17.195 136.415 17.425 ;
      RECT 137.06 19.915 137.35 20.145 ;
      RECT 135.49 19.915 135.78 20.145 ;
      RECT 133.39 19.915 133.68 20.145 ;
      RECT 133.39 19.96 137.35 20.1 ;
      RECT 137.03 22.62 137.35 22.88 ;
      RECT 136.05 22.635 136.34 22.865 ;
      RECT 136.05 22.68 137.35 22.82 ;
      RECT 137.03 28.06 137.35 28.32 ;
      RECT 136.51 28.075 136.8 28.305 ;
      RECT 136.51 28.12 137.35 28.26 ;
      RECT 136.51 16.855 136.8 17.085 ;
      RECT 136.2 16.9 136.8 17.04 ;
      RECT 136.2 16.56 136.34 17.04 ;
      RECT 134.27 16.5 134.59 16.76 ;
      RECT 134.27 16.56 136.34 16.7 ;
      RECT 131.6 17.24 135.65 17.38 ;
      RECT 135.51 16.855 135.65 17.38 ;
      RECT 131.6 16.84 131.74 17.38 ;
      RECT 131.51 16.84 131.83 17.1 ;
      RECT 135.435 16.855 135.725 17.085 ;
      RECT 134.27 27.38 134.59 27.64 ;
      RECT 135.205 27.395 135.495 27.625 ;
      RECT 134.27 27.44 135.495 27.58 ;
      RECT 134.745 16.855 135.035 17.085 ;
      RECT 132.52 16.9 135.035 17.04 ;
      RECT 132.52 16.39 132.66 17.04 ;
      RECT 129.76 16.39 132.66 16.53 ;
      RECT 128.75 16.16 129.07 16.42 ;
      RECT 129.76 16.22 129.9 16.53 ;
      RECT 128.75 16.22 129.9 16.36 ;
      RECT 134.27 22.96 134.59 23.22 ;
      RECT 131.14 23.02 134.96 23.16 ;
      RECT 134.82 22.295 134.96 23.16 ;
      RECT 131.14 22.34 131.28 23.16 ;
      RECT 128.75 22.28 129.07 22.54 ;
      RECT 123.23 22.28 123.55 22.54 ;
      RECT 117.71 22.28 118.03 22.54 ;
      RECT 134.745 22.295 135.035 22.525 ;
      RECT 124.625 22.295 124.915 22.525 ;
      RECT 110.365 22.295 110.655 22.525 ;
      RECT 110.365 22.34 131.28 22.48 ;
      RECT 134.27 14.8 134.59 15.06 ;
      RECT 133.9 14.86 134.59 15 ;
      RECT 133.9 13.795 134.04 15 ;
      RECT 133.825 13.795 134.115 14.025 ;
      RECT 134.21 19.235 134.5 19.465 ;
      RECT 134.285 18.94 134.425 19.465 ;
      RECT 131.51 18.88 131.83 19.14 ;
      RECT 131.51 18.94 134.425 19.08 ;
      RECT 128.75 19.9 129.07 20.16 ;
      RECT 128.75 19.96 131.28 20.1 ;
      RECT 131.14 19.62 131.28 20.1 ;
      RECT 132.905 19.575 133.195 19.805 ;
      RECT 131.14 19.62 133.195 19.76 ;
      RECT 121.02 14.35 128.06 14.49 ;
      RECT 127.92 14.18 128.06 14.49 ;
      RECT 131.51 14.12 131.83 14.38 ;
      RECT 121.02 14.18 121.16 14.49 ;
      RECT 127.92 14.18 131.83 14.32 ;
      RECT 120.1 14.18 121.16 14.32 ;
      RECT 120.1 13.84 120.24 14.32 ;
      RECT 118.925 13.795 119.215 14.025 ;
      RECT 118.925 13.84 120.24 13.98 ;
      RECT 131.51 17.52 131.83 17.78 ;
      RECT 128.765 17.535 129.055 17.765 ;
      RECT 128.765 17.58 131.83 17.72 ;
      RECT 131.51 21.26 131.83 21.52 ;
      RECT 125.99 21.26 126.31 21.52 ;
      RECT 125.99 21.32 131.83 21.46 ;
      RECT 127 28.12 129.9 28.26 ;
      RECT 129.76 27.78 129.9 28.26 ;
      RECT 127 27.78 127.14 28.26 ;
      RECT 131.51 27.72 131.83 27.98 ;
      RECT 120.945 27.735 121.235 27.965 ;
      RECT 129.76 27.78 131.83 27.92 ;
      RECT 122.86 27.78 127.14 27.92 ;
      RECT 122.86 27.44 123 27.92 ;
      RECT 121.02 27.44 121.16 27.965 ;
      RECT 121.02 27.44 123 27.58 ;
      RECT 125.99 26.7 126.31 26.96 ;
      RECT 131.525 26.715 131.815 26.945 ;
      RECT 125.99 26.76 131.815 26.9 ;
      RECT 129.215 21.955 129.505 22.185 ;
      RECT 126.695 21.955 126.985 22.185 ;
      RECT 125.505 21.955 125.795 22.185 ;
      RECT 125.505 22 129.505 22.14 ;
      RECT 129.215 27.395 129.505 27.625 ;
      RECT 126.695 27.395 126.985 27.625 ;
      RECT 125.505 27.395 125.795 27.625 ;
      RECT 125.505 27.44 129.505 27.58 ;
      RECT 128.75 13.78 129.07 14.04 ;
      RECT 120.765 13.795 121.055 14.025 ;
      RECT 120.765 13.84 129.07 13.98 ;
      RECT 123.23 14.8 123.55 15.06 ;
      RECT 123.23 14.86 128.98 15 ;
      RECT 128.84 14.46 128.98 15 ;
      RECT 128.75 14.46 129.07 14.72 ;
      RECT 128.75 16.84 129.07 17.1 ;
      RECT 128.075 16.855 128.365 17.085 ;
      RECT 128.075 16.9 129.07 17.04 ;
      RECT 128.75 19.22 129.07 19.48 ;
      RECT 123.23 19.22 123.55 19.48 ;
      RECT 118.72 19.28 129.07 19.42 ;
      RECT 118.72 18.94 118.86 19.42 ;
      RECT 117.71 18.88 118.03 19.14 ;
      RECT 117.71 18.94 118.86 19.08 ;
      RECT 128.78 21.615 129.07 21.845 ;
      RECT 127.21 21.615 127.5 21.845 ;
      RECT 125.11 21.615 125.4 21.845 ;
      RECT 125.11 21.66 129.07 21.8 ;
      RECT 128.78 27.055 129.07 27.285 ;
      RECT 127.21 27.055 127.5 27.285 ;
      RECT 125.11 27.055 125.4 27.285 ;
      RECT 125.11 27.1 129.07 27.24 ;
      RECT 123.23 17.18 123.55 17.44 ;
      RECT 126.925 17.195 127.215 17.425 ;
      RECT 123.23 17.24 127.215 17.38 ;
      RECT 125.99 16.84 126.31 17.1 ;
      RECT 125.99 16.855 126.435 17.085 ;
      RECT 125.99 11.4 126.31 11.66 ;
      RECT 122.785 11.415 123.075 11.645 ;
      RECT 122.785 11.46 126.31 11.6 ;
      RECT 125.99 17.52 126.31 17.78 ;
      RECT 122.4 17.58 126.31 17.72 ;
      RECT 122.4 16.855 122.54 17.72 ;
      RECT 113.125 17.195 113.415 17.425 ;
      RECT 113.125 17.24 118.4 17.38 ;
      RECT 118.26 17.07 118.4 17.38 ;
      RECT 118.26 17.07 121.62 17.21 ;
      RECT 121.48 16.9 121.62 17.21 ;
      RECT 122.325 16.855 122.615 17.085 ;
      RECT 121.48 16.9 122.615 17.04 ;
      RECT 125.99 22.62 126.31 22.88 ;
      RECT 125.93 22.635 126.31 22.865 ;
      RECT 117.34 25.06 118.86 25.2 ;
      RECT 118.72 24.72 118.86 25.2 ;
      RECT 117.34 24.38 117.48 25.2 ;
      RECT 125.99 24.66 126.31 24.92 ;
      RECT 123.32 24.72 126.31 24.86 ;
      RECT 118.72 24.72 120.7 24.86 ;
      RECT 120.56 24.38 120.7 24.86 ;
      RECT 123.32 24.38 123.46 24.86 ;
      RECT 114.045 24.335 114.335 24.565 ;
      RECT 120.56 24.38 123.46 24.52 ;
      RECT 114.045 24.38 117.48 24.52 ;
      RECT 125.99 29.42 126.31 29.68 ;
      RECT 122.785 29.435 123.075 29.665 ;
      RECT 122.785 29.48 126.31 29.62 ;
      RECT 122.785 28.415 123.075 28.645 ;
      RECT 122.785 28.46 125.3 28.6 ;
      RECT 125.16 28.12 125.3 28.6 ;
      RECT 125.93 28.075 126.22 28.305 ;
      RECT 125.16 28.12 126.22 28.26 ;
      RECT 125.545 16.855 125.835 17.085 ;
      RECT 123.32 16.9 125.835 17.04 ;
      RECT 123.32 16.16 123.46 17.04 ;
      RECT 123.23 16.16 123.55 16.42 ;
      RECT 118.11 16.16 118.43 16.42 ;
      RECT 118.11 16.22 123.55 16.36 ;
      RECT 123.23 18.54 123.55 18.8 ;
      RECT 114.95 18.54 115.27 18.8 ;
      RECT 125.085 18.555 125.375 18.785 ;
      RECT 114.95 18.6 125.375 18.74 ;
      RECT 117.71 25.68 118.03 25.94 ;
      RECT 125.085 25.695 125.375 25.925 ;
      RECT 117.71 25.74 125.375 25.88 ;
      RECT 123.23 27.38 123.55 27.64 ;
      RECT 124.625 27.395 124.915 27.625 ;
      RECT 123.23 27.44 124.915 27.58 ;
      RECT 123.23 12.08 123.55 12.34 ;
      RECT 117.71 12.08 118.03 12.34 ;
      RECT 117.71 12.14 123.55 12.28 ;
      RECT 123.23 28.06 123.55 28.32 ;
      RECT 122.17 28.12 123.55 28.26 ;
      RECT 122.17 27.735 122.31 28.26 ;
      RECT 122.095 27.735 122.385 27.965 ;
      RECT 123.23 30.1 123.55 30.36 ;
      RECT 122.095 30.115 122.385 30.345 ;
      RECT 122.095 30.16 123.55 30.3 ;
      RECT 113.2 32.88 118.86 33.02 ;
      RECT 118.72 32.2 118.86 33.02 ;
      RECT 113.2 32.2 113.34 33.02 ;
      RECT 123.23 32.14 123.55 32.4 ;
      RECT 112.19 32.14 112.51 32.4 ;
      RECT 119.49 32.155 119.78 32.385 ;
      RECT 118.72 32.2 123.55 32.34 ;
      RECT 112.19 32.2 113.34 32.34 ;
      RECT 122.775 19.575 123.065 19.805 ;
      RECT 120.255 19.575 120.545 19.805 ;
      RECT 119.065 19.575 119.355 19.805 ;
      RECT 119.065 19.62 123.065 19.76 ;
      RECT 122.775 25.015 123.065 25.245 ;
      RECT 120.255 25.015 120.545 25.245 ;
      RECT 119.065 25.015 119.355 25.245 ;
      RECT 119.065 25.06 123.065 25.2 ;
      RECT 122.34 19.915 122.63 20.145 ;
      RECT 120.77 19.915 121.06 20.145 ;
      RECT 118.67 19.915 118.96 20.145 ;
      RECT 118.67 19.96 122.63 20.1 ;
      RECT 122.34 25.355 122.63 25.585 ;
      RECT 120.77 25.355 121.06 25.585 ;
      RECT 118.67 25.355 118.96 25.585 ;
      RECT 118.67 25.4 122.63 25.54 ;
      RECT 120.47 13.1 120.79 13.36 ;
      RECT 121.405 13.115 121.695 13.345 ;
      RECT 120.47 13.16 121.695 13.3 ;
      RECT 117.71 28.06 118.03 28.32 ;
      RECT 121.405 28.075 121.695 28.305 ;
      RECT 117.71 28.12 121.695 28.26 ;
      RECT 120.945 29.775 121.235 30.005 ;
      RECT 110.44 29.65 114.26 29.79 ;
      RECT 114.12 29.48 114.26 29.79 ;
      RECT 121.02 29.48 121.16 30.005 ;
      RECT 114.95 29.42 115.27 29.68 ;
      RECT 109.43 29.42 109.75 29.68 ;
      RECT 110.44 29.48 110.58 29.79 ;
      RECT 114.12 29.48 121.16 29.62 ;
      RECT 109.43 29.48 110.58 29.62 ;
      RECT 120.47 18.88 120.79 19.14 ;
      RECT 119.49 18.895 119.78 19.125 ;
      RECT 119.49 18.94 120.79 19.08 ;
      RECT 120.47 27.04 120.79 27.3 ;
      RECT 112.19 27.04 112.51 27.3 ;
      RECT 112.19 27.1 120.79 27.24 ;
      RECT 120.47 27.72 120.79 27.98 ;
      RECT 120.255 27.735 120.79 27.965 ;
      RECT 112.19 27.72 112.51 27.98 ;
      RECT 109.43 27.72 109.75 27.98 ;
      RECT 92.87 27.72 93.19 27.98 ;
      RECT 119.565 27.735 119.855 27.965 ;
      RECT 98.94 27.78 119.855 27.92 ;
      RECT 92.87 27.78 94.02 27.92 ;
      RECT 93.88 27.44 94.02 27.92 ;
      RECT 98.94 27.44 99.08 27.92 ;
      RECT 93.88 27.44 99.08 27.58 ;
      RECT 113.2 30.5 118.86 30.64 ;
      RECT 118.72 30.16 118.86 30.64 ;
      RECT 113.2 30.16 113.34 30.64 ;
      RECT 112.19 30.1 112.51 30.36 ;
      RECT 119.565 30.115 119.855 30.345 ;
      RECT 118.72 30.16 119.855 30.3 ;
      RECT 112.19 30.16 113.34 30.3 ;
      RECT 119.49 13.455 119.78 13.685 ;
      RECT 118.26 13.5 119.78 13.64 ;
      RECT 118.26 13.33 118.4 13.64 ;
      RECT 99.4 13.33 118.4 13.47 ;
      RECT 98.39 13.1 98.71 13.36 ;
      RECT 99.4 13.16 99.54 13.47 ;
      RECT 98.39 13.16 99.54 13.3 ;
      RECT 119.49 24.335 119.78 24.565 ;
      RECT 118.72 24.38 119.78 24.52 ;
      RECT 118.72 24.04 118.86 24.52 ;
      RECT 115.885 23.995 116.175 24.225 ;
      RECT 115.885 24.04 118.86 24.18 ;
      RECT 113.2 14.69 115.64 14.83 ;
      RECT 115.5 14.52 115.64 14.83 ;
      RECT 118.11 14.46 118.43 14.72 ;
      RECT 109.43 14.46 109.75 14.72 ;
      RECT 113.2 14.52 113.34 14.83 ;
      RECT 115.5 14.52 118.43 14.66 ;
      RECT 109.43 14.52 113.34 14.66 ;
      RECT 117.8 14.18 117.94 14.66 ;
      RECT 117.8 14.18 118.4 14.32 ;
      RECT 118.26 13.795 118.4 14.32 ;
      RECT 118.185 13.795 118.475 14.025 ;
      RECT 117.71 19.56 118.03 19.82 ;
      RECT 118.185 19.575 118.475 19.805 ;
      RECT 117.71 19.62 118.475 19.76 ;
      RECT 117.71 24.66 118.03 24.92 ;
      RECT 118.185 24.675 118.475 24.905 ;
      RECT 117.71 24.72 118.475 24.86 ;
      RECT 117.71 13.78 118.03 14.04 ;
      RECT 115.425 13.795 115.715 14.025 ;
      RECT 115.425 13.84 118.03 13.98 ;
      RECT 117.71 16.84 118.03 17.1 ;
      RECT 113.815 16.855 114.105 17.085 ;
      RECT 113.815 16.9 118.03 17.04 ;
      RECT 117.71 38.26 118.03 38.52 ;
      RECT 40.43 38.26 40.75 38.52 ;
      RECT 40.43 38.32 118.03 38.46 ;
      RECT 114.95 21.26 115.27 21.52 ;
      RECT 117.265 21.275 117.555 21.505 ;
      RECT 114.95 21.32 117.555 21.46 ;
      RECT 112.19 25.68 112.51 25.94 ;
      RECT 112.19 25.74 115.41 25.88 ;
      RECT 115.27 24.675 115.41 25.88 ;
      RECT 115.195 24.675 115.485 24.905 ;
      RECT 114.95 19.22 115.27 19.48 ;
      RECT 114.505 19.235 114.795 19.465 ;
      RECT 114.505 19.28 115.27 19.42 ;
      RECT 114.955 21.955 115.245 22.185 ;
      RECT 112.435 21.955 112.725 22.185 ;
      RECT 111.245 21.955 111.535 22.185 ;
      RECT 111.245 22 115.245 22.14 ;
      RECT 114.52 21.615 114.81 21.845 ;
      RECT 112.95 21.615 113.24 21.845 ;
      RECT 110.85 21.615 111.14 21.845 ;
      RECT 110.85 21.66 114.81 21.8 ;
      RECT 112.19 17.52 112.51 17.78 ;
      RECT 114.505 17.535 114.795 17.765 ;
      RECT 112.19 17.58 114.795 17.72 ;
      RECT 109.06 25.4 111.5 25.54 ;
      RECT 111.36 25.06 111.5 25.54 ;
      RECT 109.06 25.06 109.2 25.54 ;
      RECT 111.36 25.06 114.26 25.2 ;
      RECT 114.12 24.72 114.26 25.2 ;
      RECT 96.18 25.06 109.2 25.2 ;
      RECT 82.84 25.06 85.28 25.2 ;
      RECT 85.14 24.72 85.28 25.2 ;
      RECT 66.74 25.06 72.86 25.2 ;
      RECT 72.72 24.72 72.86 25.2 ;
      RECT 57.54 25.06 61.82 25.2 ;
      RECT 61.68 24.72 61.82 25.2 ;
      RECT 96.18 24.72 96.32 25.2 ;
      RECT 82.84 24.72 82.98 25.2 ;
      RECT 66.74 24.38 66.88 25.2 ;
      RECT 57.54 24.72 57.68 25.2 ;
      RECT 114.505 24.675 114.795 24.905 ;
      RECT 22.045 24.675 22.335 24.905 ;
      RECT 114.12 24.72 114.795 24.86 ;
      RECT 92.04 24.72 96.32 24.86 ;
      RECT 85.14 24.72 89.42 24.86 ;
      RECT 89.28 24.38 89.42 24.86 ;
      RECT 72.72 24.72 82.98 24.86 ;
      RECT 61.68 24.72 65.5 24.86 ;
      RECT 65.36 24.38 65.5 24.86 ;
      RECT 56.62 24.72 57.68 24.86 ;
      RECT 23.96 24.72 45.26 24.86 ;
      RECT 45.12 24.38 45.26 24.86 ;
      RECT 92.04 24.38 92.18 24.86 ;
      RECT 56.62 23.995 56.76 24.86 ;
      RECT 23.96 24.38 24.1 24.86 ;
      RECT 22.12 24.38 22.26 24.905 ;
      RECT 45.95 24.32 46.27 24.58 ;
      RECT 89.28 24.38 92.18 24.52 ;
      RECT 65.36 24.38 66.88 24.52 ;
      RECT 52.48 24.38 55.84 24.52 ;
      RECT 55.7 24.04 55.84 24.52 ;
      RECT 45.12 24.38 49.4 24.52 ;
      RECT 49.26 24.04 49.4 24.52 ;
      RECT 22.12 24.38 24.1 24.52 ;
      RECT 52.48 24.04 52.62 24.52 ;
      RECT 56.545 23.995 56.835 24.225 ;
      RECT 55.7 24.04 56.835 24.18 ;
      RECT 49.26 24.04 52.62 24.18 ;
      RECT 113.355 24.675 113.645 24.905 ;
      RECT 113.43 24.04 113.57 24.905 ;
      RECT 112.19 23.98 112.51 24.24 ;
      RECT 112.19 24.04 113.57 24.18 ;
      RECT 97.025 17.24 98.62 17.38 ;
      RECT 98.48 16.9 98.62 17.38 ;
      RECT 97.025 16.9 97.165 17.38 ;
      RECT 101.15 16.84 101.47 17.1 ;
      RECT 112.665 16.855 112.955 17.085 ;
      RECT 103.465 16.855 103.755 17.085 ;
      RECT 96.105 16.855 96.395 17.085 ;
      RECT 108.6 16.9 109.66 17.04 ;
      RECT 109.52 16.56 109.66 17.04 ;
      RECT 98.48 16.9 106.44 17.04 ;
      RECT 106.3 16.56 106.44 17.04 ;
      RECT 96.105 16.9 97.165 17.04 ;
      RECT 108.6 16.56 108.74 17.04 ;
      RECT 112.74 16.56 112.88 17.085 ;
      RECT 109.52 16.56 112.88 16.7 ;
      RECT 106.3 16.56 108.74 16.7 ;
      RECT 109.43 24.66 109.75 24.92 ;
      RECT 112.665 24.675 112.955 24.905 ;
      RECT 109.43 24.72 112.955 24.86 ;
      RECT 98.02 14.18 102.76 14.32 ;
      RECT 102.62 13.84 102.76 14.32 ;
      RECT 98.02 13.5 98.16 14.32 ;
      RECT 112.19 13.78 112.51 14.04 ;
      RECT 103.465 13.795 103.755 14.025 ;
      RECT 102.62 13.84 112.51 13.98 ;
      RECT 94.725 13.455 95.015 13.685 ;
      RECT 94.725 13.5 98.16 13.64 ;
      RECT 112.19 15.82 112.51 16.08 ;
      RECT 109.43 15.82 109.75 16.08 ;
      RECT 109.43 15.88 112.51 16.02 ;
      RECT 112.19 16.84 112.51 17.1 ;
      RECT 111.975 16.855 112.51 17.085 ;
      RECT 112.19 22.62 112.51 22.88 ;
      RECT 111.67 22.635 111.96 22.865 ;
      RECT 111.67 22.68 112.51 22.82 ;
      RECT 87.35 31.12 87.67 31.38 ;
      RECT 76.31 31.12 76.63 31.38 ;
      RECT 80.54 31.18 88.5 31.32 ;
      RECT 88.36 31.01 88.5 31.32 ;
      RECT 76.31 31.18 77.46 31.32 ;
      RECT 77.32 30.84 77.46 31.32 ;
      RECT 83.76 30.16 83.9 31.32 ;
      RECT 80.54 30.84 80.68 31.32 ;
      RECT 88.36 31.01 96.55 31.15 ;
      RECT 96.41 30.115 96.55 31.15 ;
      RECT 112.19 30.78 112.51 31.04 ;
      RECT 111.36 30.84 112.51 30.98 ;
      RECT 96.41 30.84 101.38 30.98 ;
      RECT 101.24 30.5 101.38 30.98 ;
      RECT 77.32 30.84 80.68 30.98 ;
      RECT 111.36 30.5 111.5 30.98 ;
      RECT 101.24 30.5 111.5 30.64 ;
      RECT 96.335 30.115 96.625 30.345 ;
      RECT 82.995 30.115 83.285 30.345 ;
      RECT 82.995 30.16 83.9 30.3 ;
      RECT 109.43 17.52 109.75 17.78 ;
      RECT 103.91 17.52 104.23 17.78 ;
      RECT 108.6 17.58 111.5 17.72 ;
      RECT 111.36 16.855 111.5 17.72 ;
      RECT 103.91 17.58 105.06 17.72 ;
      RECT 104.92 17.41 105.06 17.72 ;
      RECT 108.6 17.41 108.74 17.72 ;
      RECT 104.92 17.41 108.74 17.55 ;
      RECT 111.285 16.855 111.575 17.085 ;
      RECT 97.945 16.855 98.235 17.085 ;
      RECT 98.02 15.88 98.16 17.085 ;
      RECT 88.82 16.05 97.24 16.19 ;
      RECT 97.1 15.88 97.24 16.19 ;
      RECT 103.91 15.82 104.23 16.08 ;
      RECT 87.35 15.82 87.67 16.08 ;
      RECT 88.82 15.88 88.96 16.19 ;
      RECT 97.1 15.88 104.23 16.02 ;
      RECT 87.35 15.88 88.96 16.02 ;
      RECT 101.15 21.26 101.47 21.52 ;
      RECT 102.545 21.275 102.835 21.505 ;
      RECT 101.15 21.32 102.835 21.46 ;
      RECT 101.15 22.62 101.47 22.88 ;
      RECT 96.95 22.635 97.24 22.865 ;
      RECT 96.95 22.68 101.47 22.82 ;
      RECT 98.02 29.82 100.46 29.96 ;
      RECT 100.32 29.48 100.46 29.96 ;
      RECT 98.02 29.48 98.16 29.96 ;
      RECT 101.15 29.42 101.47 29.68 ;
      RECT 97.025 29.435 97.315 29.665 ;
      RECT 100.32 29.48 101.47 29.62 ;
      RECT 97.025 29.48 98.16 29.62 ;
      RECT 96.64 18.94 100 19.08 ;
      RECT 99.86 18.6 100 19.08 ;
      RECT 96.64 18.6 96.78 19.08 ;
      RECT 87.35 18.54 87.67 18.8 ;
      RECT 100.705 18.555 100.995 18.785 ;
      RECT 99.86 18.6 100.995 18.74 ;
      RECT 87.35 18.6 96.78 18.74 ;
      RECT 95.63 20.24 95.95 20.5 ;
      RECT 100.705 20.255 100.995 20.485 ;
      RECT 95.63 20.3 100.995 20.44 ;
      RECT 100.235 21.955 100.525 22.185 ;
      RECT 97.715 21.955 98.005 22.185 ;
      RECT 96.525 21.955 96.815 22.185 ;
      RECT 96.525 22 100.525 22.14 ;
      RECT 99.8 21.615 100.09 21.845 ;
      RECT 98.23 21.615 98.52 21.845 ;
      RECT 96.13 21.615 96.42 21.845 ;
      RECT 96.13 21.66 100.09 21.8 ;
      RECT 98.39 23.98 98.71 24.24 ;
      RECT 97.945 23.995 98.235 24.225 ;
      RECT 97.945 24.04 98.71 24.18 ;
      RECT 90.11 28.4 90.43 28.66 ;
      RECT 97.56 28.46 98.62 28.6 ;
      RECT 98.48 28.06 98.62 28.6 ;
      RECT 90.11 28.46 91.26 28.6 ;
      RECT 91.12 28.29 91.26 28.6 ;
      RECT 97.56 28.29 97.7 28.6 ;
      RECT 91.12 28.29 97.7 28.43 ;
      RECT 98.39 28.06 98.71 28.32 ;
      RECT 98.395 19.575 98.685 19.805 ;
      RECT 95.875 19.575 96.165 19.805 ;
      RECT 94.685 19.575 94.975 19.805 ;
      RECT 94.685 19.62 98.685 19.76 ;
      RECT 97.96 19.915 98.25 20.145 ;
      RECT 96.39 19.915 96.68 20.145 ;
      RECT 94.29 19.915 94.58 20.145 ;
      RECT 94.29 19.96 98.25 20.1 ;
      RECT 97.34 16.855 97.63 17.085 ;
      RECT 83.915 16.855 84.205 17.085 ;
      RECT 97.415 16.56 97.555 17.085 ;
      RECT 83.99 16.22 84.13 17.085 ;
      RECT 92.87 16.5 93.19 16.76 ;
      RECT 87.9 16.56 97.555 16.7 ;
      RECT 87.9 16.22 88.04 16.7 ;
      RECT 84.59 16.16 84.91 16.42 ;
      RECT 83.99 16.22 88.04 16.36 ;
      RECT 81.83 17.52 82.15 17.78 ;
      RECT 73.55 17.52 73.87 17.78 ;
      RECT 73.55 17.58 75.16 17.72 ;
      RECT 75.02 17.41 75.16 17.72 ;
      RECT 74.1 16.855 74.24 17.72 ;
      RECT 82.84 17.41 88.04 17.55 ;
      RECT 87.9 17.24 88.04 17.55 ;
      RECT 75.02 17.41 78.84 17.55 ;
      RECT 78.7 17.24 78.84 17.55 ;
      RECT 81.92 17.24 82.06 17.78 ;
      RECT 96.565 17.195 96.855 17.425 ;
      RECT 82.84 17.24 82.98 17.55 ;
      RECT 87.9 17.24 96.855 17.38 ;
      RECT 78.7 17.24 82.98 17.38 ;
      RECT 74.025 16.855 74.315 17.085 ;
      RECT 95.63 13.1 95.95 13.36 ;
      RECT 96.1 13.115 96.39 13.345 ;
      RECT 95.63 13.16 96.39 13.3 ;
      RECT 95.63 13.78 95.95 14.04 ;
      RECT 95.415 13.795 95.95 14.025 ;
      RECT 95.63 16.84 95.95 17.1 ;
      RECT 95.415 16.855 95.95 17.085 ;
      RECT 87.35 19.56 87.67 19.82 ;
      RECT 85.37 19.62 92.64 19.76 ;
      RECT 92.5 19.28 92.64 19.76 ;
      RECT 85.37 19.235 85.51 19.76 ;
      RECT 85.295 19.235 85.585 19.465 ;
      RECT 92.5 19.28 95.86 19.42 ;
      RECT 95.72 18.88 95.86 19.42 ;
      RECT 95.63 18.88 95.95 19.14 ;
      RECT 92.35 24.335 92.64 24.565 ;
      RECT 92.425 24.04 92.565 24.565 ;
      RECT 95.63 23.98 95.95 24.24 ;
      RECT 92.425 24.04 95.95 24.18 ;
      RECT 95.185 29.775 95.475 30.005 ;
      RECT 95.185 29.82 95.86 29.96 ;
      RECT 95.72 29.42 95.86 29.96 ;
      RECT 95.63 29.42 95.95 29.68 ;
      RECT 81.83 22.96 82.15 23.22 ;
      RECT 80.465 22.975 80.755 23.205 ;
      RECT 80.465 23.02 82.15 23.16 ;
      RECT 81 22.295 81.14 23.16 ;
      RECT 92.87 22.28 93.19 22.54 ;
      RECT 90.11 22.28 90.43 22.54 ;
      RECT 95.645 22.295 95.935 22.525 ;
      RECT 80.925 22.295 81.215 22.525 ;
      RECT 80.925 22.34 95.935 22.48 ;
      RECT 95.635 25.015 95.925 25.245 ;
      RECT 93.115 25.015 93.405 25.245 ;
      RECT 91.925 25.015 92.215 25.245 ;
      RECT 91.925 25.06 95.925 25.2 ;
      RECT 95.2 25.355 95.49 25.585 ;
      RECT 93.63 25.355 93.92 25.585 ;
      RECT 91.53 25.355 91.82 25.585 ;
      RECT 91.53 25.4 95.49 25.54 ;
      RECT 92.87 18.88 93.19 19.14 ;
      RECT 95.11 18.895 95.4 19.125 ;
      RECT 92.87 18.94 95.4 19.08 ;
      RECT 92.87 17.52 93.19 17.78 ;
      RECT 94.725 17.535 95.015 17.765 ;
      RECT 92.87 17.58 95.015 17.72 ;
      RECT 84.59 30.44 84.91 30.7 ;
      RECT 84.59 30.5 94.71 30.64 ;
      RECT 94.57 30.115 94.71 30.64 ;
      RECT 94.495 30.115 94.785 30.345 ;
      RECT 90.11 14.46 90.43 14.72 ;
      RECT 90.11 14.52 94.48 14.66 ;
      RECT 94.34 13.795 94.48 14.66 ;
      RECT 94.265 13.795 94.555 14.025 ;
      RECT 92.87 19.56 93.19 19.82 ;
      RECT 93.805 19.575 94.095 19.805 ;
      RECT 92.87 19.62 94.095 19.76 ;
      RECT 93.805 30.115 94.095 30.345 ;
      RECT 93.88 29.82 94.02 30.345 ;
      RECT 92.87 29.76 93.19 30.02 ;
      RECT 92.87 29.82 94.02 29.96 ;
      RECT 93.575 13.795 93.865 14.025 ;
      RECT 93.65 13.16 93.79 14.025 ;
      RECT 92.87 13.1 93.19 13.36 ;
      RECT 92.87 13.16 93.79 13.3 ;
      RECT 92.87 22.96 93.19 23.22 ;
      RECT 82.335 23.02 93.19 23.16 ;
      RECT 82.335 22.635 82.475 23.16 ;
      RECT 82.26 22.635 82.55 22.865 ;
      RECT 84.59 27.38 84.91 27.64 ;
      RECT 84.59 27.44 92.18 27.58 ;
      RECT 92.04 27.1 92.18 27.58 ;
      RECT 92.87 27.04 93.19 27.3 ;
      RECT 92.04 27.1 93.19 27.24 ;
      RECT 87.35 14.8 87.67 15.06 ;
      RECT 87.44 13.84 87.58 15.06 ;
      RECT 71.8 14.18 74.24 14.32 ;
      RECT 74.1 13.84 74.24 14.32 ;
      RECT 71.8 13.84 71.94 14.32 ;
      RECT 82.215 13.78 82.535 14.04 ;
      RECT 70.79 13.78 71.11 14.04 ;
      RECT 92.885 13.795 93.175 14.025 ;
      RECT 63.905 13.795 64.195 14.025 ;
      RECT 74.1 13.84 93.175 13.98 ;
      RECT 69.04 13.84 71.94 13.98 ;
      RECT 63.905 13.84 66.42 13.98 ;
      RECT 66.28 13.5 66.42 13.98 ;
      RECT 69.04 13.5 69.18 13.98 ;
      RECT 66.28 13.5 69.18 13.64 ;
      RECT 90.11 11.4 90.43 11.66 ;
      RECT 91.505 11.415 91.795 11.645 ;
      RECT 90.11 11.46 91.795 11.6 ;
      RECT 90.11 24.66 90.43 24.92 ;
      RECT 91.045 24.675 91.335 24.905 ;
      RECT 90.11 24.72 91.335 24.86 ;
      RECT 84.605 19.235 84.895 19.465 ;
      RECT 86.98 19.11 89.42 19.25 ;
      RECT 89.28 18.94 89.42 19.25 ;
      RECT 84.68 18.94 84.82 19.465 ;
      RECT 90.11 18.88 90.43 19.14 ;
      RECT 86.98 18.94 87.12 19.25 ;
      RECT 89.28 18.94 90.43 19.08 ;
      RECT 84.68 18.94 87.12 19.08 ;
      RECT 90.11 21.26 90.43 21.52 ;
      RECT 87.825 21.275 88.115 21.505 ;
      RECT 87.825 21.32 90.43 21.46 ;
      RECT 90.11 29.76 90.43 30.02 ;
      RECT 82.345 29.775 82.635 30.005 ;
      RECT 82.345 29.82 90.43 29.96 ;
      RECT 87.35 11.74 87.67 12 ;
      RECT 87.44 11.46 87.58 12 ;
      RECT 81.83 11.4 82.15 11.66 ;
      RECT 82.765 11.415 83.055 11.645 ;
      RECT 81.83 11.46 87.58 11.6 ;
      RECT 87.35 16.84 87.67 17.1 ;
      RECT 84.605 16.855 84.895 17.085 ;
      RECT 84.605 16.9 87.67 17.04 ;
      RECT 84.59 20.24 84.91 20.5 ;
      RECT 85.985 20.255 86.275 20.485 ;
      RECT 84.59 20.3 86.275 20.44 ;
      RECT 85.515 21.955 85.805 22.185 ;
      RECT 82.995 21.955 83.285 22.185 ;
      RECT 81.805 21.955 82.095 22.185 ;
      RECT 81.805 22 85.805 22.14 ;
      RECT 85.08 21.615 85.37 21.845 ;
      RECT 83.51 21.615 83.8 21.845 ;
      RECT 81.41 21.615 81.7 21.845 ;
      RECT 81.41 21.66 85.37 21.8 ;
      RECT 84.145 18.895 84.435 19.125 ;
      RECT 84.22 18.6 84.36 19.125 ;
      RECT 84.59 18.54 84.91 18.8 ;
      RECT 84.22 18.6 84.91 18.74 ;
      RECT 67.51 22.295 67.8 22.525 ;
      RECT 67.51 22.34 71.94 22.48 ;
      RECT 71.8 22 71.94 22.48 ;
      RECT 71.8 22 74.7 22.14 ;
      RECT 74.56 21.66 74.7 22.14 ;
      RECT 74.56 21.66 81.14 21.8 ;
      RECT 81 21.32 81.14 21.8 ;
      RECT 84.59 21.26 84.91 21.52 ;
      RECT 81 21.32 84.91 21.46 ;
      RECT 80.08 24.21 83.44 24.35 ;
      RECT 83.3 24.04 83.44 24.35 ;
      RECT 70.88 24.21 77.92 24.35 ;
      RECT 77.78 24.04 77.92 24.35 ;
      RECT 84.59 23.98 84.91 24.24 ;
      RECT 68.03 23.98 68.35 24.24 ;
      RECT 84.145 23.995 84.435 24.225 ;
      RECT 80.08 24.04 80.22 24.35 ;
      RECT 70.88 24.04 71.02 24.35 ;
      RECT 83.3 24.04 84.91 24.18 ;
      RECT 77.78 24.04 80.22 24.18 ;
      RECT 68.03 24.04 71.02 24.18 ;
      RECT 84.59 29.42 84.91 29.68 ;
      RECT 83.685 29.435 83.975 29.665 ;
      RECT 83.685 29.48 84.91 29.62 ;
      RECT 77.32 32.88 81.14 33.02 ;
      RECT 81 32.2 81.14 33.02 ;
      RECT 77.32 32.2 77.46 33.02 ;
      RECT 84.59 32.14 84.91 32.4 ;
      RECT 81.83 32.14 82.15 32.4 ;
      RECT 73.55 32.14 73.87 32.4 ;
      RECT 81 32.2 84.91 32.34 ;
      RECT 73.55 32.2 77.46 32.34 ;
      RECT 79.07 20.24 79.39 20.5 ;
      RECT 71.34 20.3 83.44 20.44 ;
      RECT 83.3 19.96 83.44 20.44 ;
      RECT 71.34 19.62 71.48 20.44 ;
      RECT 83.3 19.96 83.67 20.1 ;
      RECT 83.53 19.235 83.67 20.1 ;
      RECT 71.195 19.62 71.48 19.76 ;
      RECT 71.195 19.235 71.335 19.76 ;
      RECT 83.455 19.235 83.745 19.465 ;
      RECT 71.12 19.235 71.41 19.465 ;
      RECT 83.225 16.855 83.515 17.085 ;
      RECT 83.3 15.88 83.44 17.085 ;
      RECT 77.78 16.05 81.14 16.19 ;
      RECT 81 15.88 81.14 16.19 ;
      RECT 73.55 15.82 73.87 16.08 ;
      RECT 77.78 15.88 77.92 16.19 ;
      RECT 81 15.88 83.44 16.02 ;
      RECT 73.55 15.88 77.92 16.02 ;
      RECT 82.765 16.855 83.055 17.085 ;
      RECT 82.84 16.22 82.98 17.085 ;
      RECT 81.83 16.16 82.15 16.42 ;
      RECT 81.83 16.22 82.98 16.36 ;
      RECT 81.83 19.56 82.15 19.82 ;
      RECT 71.8 19.62 76.08 19.76 ;
      RECT 75.94 19.28 76.08 19.76 ;
      RECT 71.8 19.235 71.94 19.76 ;
      RECT 81.92 19.28 82.06 19.82 ;
      RECT 82.765 19.235 83.055 19.465 ;
      RECT 71.725 19.235 72.015 19.465 ;
      RECT 75.94 19.28 83.055 19.42 ;
      RECT 81.83 18.88 82.15 19.14 ;
      RECT 81.83 18.94 82.52 19.08 ;
      RECT 82.38 18.555 82.52 19.08 ;
      RECT 82.305 18.555 82.595 18.785 ;
      RECT 60.76 17.41 63.2 17.55 ;
      RECT 63.06 17.24 63.2 17.55 ;
      RECT 56.99 17.18 57.31 17.44 ;
      RECT 60.76 17.24 60.9 17.55 ;
      RECT 63.06 17.24 69.41 17.38 ;
      RECT 69.27 16.855 69.41 17.38 ;
      RECT 48.34 17.24 60.9 17.38 ;
      RECT 67.66 15.88 67.8 17.38 ;
      RECT 48.34 16.9 48.48 17.38 ;
      RECT 82.075 16.855 82.365 17.085 ;
      RECT 69.195 16.855 69.485 17.085 ;
      RECT 47.115 16.855 47.405 17.085 ;
      RECT 47.115 16.9 48.48 17.04 ;
      RECT 82.15 16.56 82.29 17.085 ;
      RECT 76.86 16.56 82.29 16.7 ;
      RECT 76.86 16.22 77 16.7 ;
      RECT 72.26 16.22 77 16.36 ;
      RECT 72.26 15.88 72.4 16.36 ;
      RECT 67.66 15.88 72.4 16.02 ;
      RECT 81.83 30.78 82.15 31.04 ;
      RECT 81.23 30.84 82.15 30.98 ;
      RECT 81.23 30.115 81.37 30.98 ;
      RECT 81.155 30.115 81.445 30.345 ;
      RECT 75.865 29.775 76.155 30.005 ;
      RECT 75.865 29.82 81.14 29.96 ;
      RECT 81.845 29.715 82.135 29.945 ;
      RECT 81 29.76 82.135 29.9 ;
      RECT 75.94 29.48 76.08 30.005 ;
      RECT 76.31 29.42 76.63 29.68 ;
      RECT 75.94 29.48 76.63 29.62 ;
      RECT 81.835 25.015 82.125 25.245 ;
      RECT 79.315 25.015 79.605 25.245 ;
      RECT 78.125 25.015 78.415 25.245 ;
      RECT 78.125 25.06 82.125 25.2 ;
      RECT 81.4 25.355 81.69 25.585 ;
      RECT 79.83 25.355 80.12 25.585 ;
      RECT 77.73 25.355 78.02 25.585 ;
      RECT 77.73 25.4 81.69 25.54 ;
      RECT 79.07 17.52 79.39 17.78 ;
      RECT 81.385 17.535 81.675 17.765 ;
      RECT 79.07 17.58 81.675 17.72 ;
      RECT 79.07 30.1 79.39 30.36 ;
      RECT 80.465 30.115 80.755 30.345 ;
      RECT 79.07 30.16 80.755 30.3 ;
      RECT 79.995 19.575 80.285 19.805 ;
      RECT 77.475 19.575 77.765 19.805 ;
      RECT 76.285 19.575 76.575 19.805 ;
      RECT 76.285 19.62 80.285 19.76 ;
      RECT 79.56 19.915 79.85 20.145 ;
      RECT 77.99 19.915 78.28 20.145 ;
      RECT 75.89 19.915 76.18 20.145 ;
      RECT 75.89 19.96 79.85 20.1 ;
      RECT 71.195 17.24 72.86 17.38 ;
      RECT 72.72 16.56 72.86 17.38 ;
      RECT 71.195 16.855 71.335 17.38 ;
      RECT 79.07 16.84 79.39 17.1 ;
      RECT 71.12 16.855 71.41 17.085 ;
      RECT 74.56 16.9 79.39 17.04 ;
      RECT 74.56 16.56 74.7 17.04 ;
      RECT 73.55 16.5 73.87 16.76 ;
      RECT 72.72 16.56 74.7 16.7 ;
      RECT 79.07 18.88 79.39 19.14 ;
      RECT 76.71 18.895 77 19.125 ;
      RECT 76.71 18.94 79.39 19.08 ;
      RECT 79.07 24.32 79.39 24.58 ;
      RECT 78.55 24.335 78.84 24.565 ;
      RECT 78.55 24.38 79.39 24.52 ;
      RECT 79.07 29.42 79.39 29.68 ;
      RECT 77.245 29.435 77.535 29.665 ;
      RECT 77.245 29.48 79.39 29.62 ;
      RECT 73.55 25 73.87 25.26 ;
      RECT 77.245 25.015 77.535 25.245 ;
      RECT 73.55 25.06 77.535 25.2 ;
      RECT 76.31 30.1 76.63 30.36 ;
      RECT 76.31 30.115 76.845 30.345 ;
      RECT 76.31 22.96 76.63 23.22 ;
      RECT 73.105 22.975 73.395 23.205 ;
      RECT 73.105 23.02 76.63 23.16 ;
      RECT 73.18 33.22 75.62 33.36 ;
      RECT 75.48 32.54 75.62 33.36 ;
      RECT 73.18 32.88 73.32 33.36 ;
      RECT 66.28 32.88 73.32 33.02 ;
      RECT 66.28 32.54 66.42 33.02 ;
      RECT 76.31 32.48 76.63 32.74 ;
      RECT 65.27 32.48 65.59 32.74 ;
      RECT 75.48 32.54 76.63 32.68 ;
      RECT 65.27 32.54 66.42 32.68 ;
      RECT 73.55 19.22 73.87 19.48 ;
      RECT 75.405 19.235 75.695 19.465 ;
      RECT 73.55 19.28 75.695 19.42 ;
      RECT 75.405 29.775 75.695 30.005 ;
      RECT 74.1 29.82 75.695 29.96 ;
      RECT 74.1 29.48 74.24 29.96 ;
      RECT 73.55 29.42 73.87 29.68 ;
      RECT 73.55 29.48 74.24 29.62 ;
      RECT 73.55 30.78 73.87 31.04 ;
      RECT 73.55 30.84 74.93 30.98 ;
      RECT 74.79 30.115 74.93 30.98 ;
      RECT 74.715 30.115 75.005 30.345 ;
      RECT 73.55 11.4 73.87 11.66 ;
      RECT 74.025 11.415 74.315 11.645 ;
      RECT 73.55 11.46 74.315 11.6 ;
      RECT 73.55 30.1 73.87 30.36 ;
      RECT 74.025 30.115 74.315 30.345 ;
      RECT 63.06 30.16 74.315 30.3 ;
      RECT 63.06 29.48 63.2 30.3 ;
      RECT 55.24 29.82 58.6 29.96 ;
      RECT 58.46 29.48 58.6 29.96 ;
      RECT 55.24 29.65 55.38 29.96 ;
      RECT 48.8 29.65 55.38 29.79 ;
      RECT 45.95 29.42 46.27 29.68 ;
      RECT 48.8 29.48 48.94 29.79 ;
      RECT 58.46 29.48 63.2 29.62 ;
      RECT 45.95 29.48 48.94 29.62 ;
      RECT 73.55 28.4 73.87 28.66 ;
      RECT 73.55 28.46 74.24 28.6 ;
      RECT 74.1 26.76 74.24 28.6 ;
      RECT 69.885 27.735 70.175 27.965 ;
      RECT 69.96 26.76 70.1 27.965 ;
      RECT 62.51 26.7 62.83 26.96 ;
      RECT 66.205 26.715 66.495 26.945 ;
      RECT 62.51 26.76 74.24 26.9 ;
      RECT 62.065 13.455 62.355 13.685 ;
      RECT 62.065 13.5 62.74 13.64 ;
      RECT 62.6 13.1 62.74 13.64 ;
      RECT 73.55 13.1 73.87 13.36 ;
      RECT 62.51 13.1 62.83 13.36 ;
      RECT 62.51 13.16 73.87 13.3 ;
      RECT 69.885 18.895 70.175 19.125 ;
      RECT 69.885 18.94 72.4 19.08 ;
      RECT 72.26 18.6 72.4 19.08 ;
      RECT 73.55 18.54 73.87 18.8 ;
      RECT 72.26 18.6 73.87 18.74 ;
      RECT 71.035 27.735 71.325 27.965 ;
      RECT 71.11 27.44 71.25 27.965 ;
      RECT 71.11 27.44 73.78 27.58 ;
      RECT 73.64 27.04 73.78 27.58 ;
      RECT 73.55 27.04 73.87 27.3 ;
      RECT 73.55 27.72 73.87 27.98 ;
      RECT 71.725 27.735 72.015 27.965 ;
      RECT 71.725 27.78 73.87 27.92 ;
      RECT 71.69 16.855 71.98 17.085 ;
      RECT 71.765 16.22 71.905 17.085 ;
      RECT 70.79 16.16 71.11 16.42 ;
      RECT 70.79 16.22 71.905 16.36 ;
      RECT 70.79 17.52 71.11 17.78 ;
      RECT 70.88 17.24 71.02 17.78 ;
      RECT 70.345 17.195 70.635 17.425 ;
      RECT 70.345 17.24 71.02 17.38 ;
      RECT 70.79 31.12 71.11 31.38 ;
      RECT 66.205 31.135 66.495 31.365 ;
      RECT 69.96 31.18 71.11 31.32 ;
      RECT 58.92 31.18 67.34 31.32 ;
      RECT 67.2 30.84 67.34 31.32 ;
      RECT 69.96 30.84 70.1 31.32 ;
      RECT 58.92 30.5 59.06 31.32 ;
      RECT 67.2 30.84 70.1 30.98 ;
      RECT 47.88 30.5 59.06 30.64 ;
      RECT 47.88 29.775 48.02 30.64 ;
      RECT 40.43 29.76 40.75 30.02 ;
      RECT 47.805 29.775 48.095 30.005 ;
      RECT 40.43 29.82 48.095 29.96 ;
      RECT 70.795 21.955 71.085 22.185 ;
      RECT 68.275 21.955 68.565 22.185 ;
      RECT 67.085 21.955 67.375 22.185 ;
      RECT 67.085 22 71.085 22.14 ;
      RECT 70.36 21.615 70.65 21.845 ;
      RECT 68.79 21.615 69.08 21.845 ;
      RECT 66.69 21.615 66.98 21.845 ;
      RECT 66.69 21.66 70.65 21.8 ;
      RECT 65.27 19.56 65.59 19.82 ;
      RECT 65.27 19.62 70.56 19.76 ;
      RECT 70.42 19.235 70.56 19.76 ;
      RECT 70.345 19.235 70.635 19.465 ;
      RECT 56.99 28.06 57.31 28.32 ;
      RECT 70.345 28.075 70.635 28.305 ;
      RECT 47.805 28.075 48.095 28.305 ;
      RECT 52.02 28.12 70.635 28.26 ;
      RECT 42.82 28.12 49.86 28.26 ;
      RECT 49.72 27.95 49.86 28.26 ;
      RECT 52.02 27.95 52.16 28.26 ;
      RECT 42.82 27.78 42.96 28.26 ;
      RECT 49.72 27.95 52.16 28.09 ;
      RECT 40.445 27.735 40.735 27.965 ;
      RECT 40.445 27.78 42.96 27.92 ;
      RECT 69.885 16.855 70.175 17.085 ;
      RECT 69.96 16.56 70.1 17.085 ;
      RECT 68.03 16.5 68.35 16.76 ;
      RECT 68.03 16.56 70.1 16.7 ;
      RECT 69.195 19.235 69.485 19.465 ;
      RECT 68.12 19.28 69.485 19.42 ;
      RECT 68.12 19.11 68.26 19.42 ;
      RECT 61.22 19.11 68.26 19.25 ;
      RECT 61.22 18.6 61.36 19.25 ;
      RECT 56.99 18.54 57.31 18.8 ;
      RECT 56.99 18.6 61.36 18.74 ;
      RECT 69.195 27.735 69.485 27.965 ;
      RECT 69.27 27.44 69.41 27.965 ;
      RECT 65.27 27.38 65.59 27.64 ;
      RECT 65.27 27.44 69.41 27.58 ;
      RECT 68.03 17.52 68.35 17.78 ;
      RECT 68.505 17.535 68.795 17.765 ;
      RECT 68.03 17.58 68.795 17.72 ;
      RECT 54.23 20.24 54.55 20.5 ;
      RECT 68.505 20.255 68.795 20.485 ;
      RECT 67.66 20.3 68.795 20.44 ;
      RECT 58.46 20.3 64.58 20.44 ;
      RECT 64.44 20.13 64.58 20.44 ;
      RECT 54.23 20.3 55.38 20.44 ;
      RECT 55.24 19.96 55.38 20.44 ;
      RECT 67.66 20.13 67.8 20.44 ;
      RECT 58.46 19.96 58.6 20.44 ;
      RECT 64.44 20.13 67.8 20.27 ;
      RECT 55.24 19.96 58.6 20.1 ;
      RECT 62.51 28.4 62.83 28.66 ;
      RECT 68.505 28.415 68.795 28.645 ;
      RECT 62.51 28.46 68.795 28.6 ;
      RECT 68.03 14.8 68.35 15.06 ;
      RECT 67.66 14.86 68.35 15 ;
      RECT 67.66 13.84 67.8 15 ;
      RECT 66.665 13.795 66.955 14.025 ;
      RECT 66.665 13.84 67.8 13.98 ;
      RECT 68.03 27.72 68.35 27.98 ;
      RECT 60.61 27.735 60.9 27.965 ;
      RECT 60.61 27.78 68.35 27.92 ;
      RECT 65.27 15.82 65.59 16.08 ;
      RECT 66.205 15.835 66.495 16.065 ;
      RECT 65.27 15.88 66.495 16.02 ;
      RECT 62.51 18.54 62.83 18.8 ;
      RECT 66.205 18.555 66.495 18.785 ;
      RECT 62.51 18.6 66.495 18.74 ;
      RECT 65.27 22.28 65.59 22.54 ;
      RECT 66.205 22.295 66.495 22.525 ;
      RECT 51.485 22.295 51.775 22.525 ;
      RECT 65.27 22.34 66.495 22.48 ;
      RECT 51.485 22.34 60.9 22.48 ;
      RECT 60.76 22 60.9 22.48 ;
      RECT 65.36 22 65.5 22.54 ;
      RECT 60.76 22 65.5 22.14 ;
      RECT 62.51 25.34 62.83 25.6 ;
      RECT 62.51 25.4 65.96 25.54 ;
      RECT 65.82 24.675 65.96 25.54 ;
      RECT 65.745 24.675 66.035 24.905 ;
      RECT 65.27 12.08 65.59 12.34 ;
      RECT 51.47 12.08 51.79 12.34 ;
      RECT 64.44 12.14 65.59 12.28 ;
      RECT 51.47 12.14 52.62 12.28 ;
      RECT 52.48 11.46 52.62 12.28 ;
      RECT 64.44 11.97 64.58 12.28 ;
      RECT 61.68 11.97 64.58 12.11 ;
      RECT 51.56 11.46 51.7 12.34 ;
      RECT 61.68 11.46 61.82 12.11 ;
      RECT 48.725 11.415 49.015 11.645 ;
      RECT 52.48 11.46 61.82 11.6 ;
      RECT 48.725 11.46 51.7 11.6 ;
      RECT 63.895 16.515 64.185 16.745 ;
      RECT 61.375 16.515 61.665 16.745 ;
      RECT 60.185 16.515 60.475 16.745 ;
      RECT 60.185 16.56 64.185 16.7 ;
      RECT 63.895 19.575 64.185 19.805 ;
      RECT 61.375 19.575 61.665 19.805 ;
      RECT 60.185 19.575 60.475 19.805 ;
      RECT 60.185 19.62 64.185 19.76 ;
      RECT 63.895 27.395 64.185 27.625 ;
      RECT 61.375 27.395 61.665 27.625 ;
      RECT 60.185 27.395 60.475 27.625 ;
      RECT 60.185 27.44 64.185 27.58 ;
      RECT 63.895 30.455 64.185 30.685 ;
      RECT 61.375 30.455 61.665 30.685 ;
      RECT 60.185 30.455 60.475 30.685 ;
      RECT 60.185 30.5 64.185 30.64 ;
      RECT 63.46 16.175 63.75 16.405 ;
      RECT 61.89 16.175 62.18 16.405 ;
      RECT 59.79 16.175 60.08 16.405 ;
      RECT 59.79 16.22 63.75 16.36 ;
      RECT 63.46 19.915 63.75 20.145 ;
      RECT 61.89 19.915 62.18 20.145 ;
      RECT 59.79 19.915 60.08 20.145 ;
      RECT 59.79 19.96 63.75 20.1 ;
      RECT 63.46 27.055 63.75 27.285 ;
      RECT 61.89 27.055 62.18 27.285 ;
      RECT 59.79 27.055 60.08 27.285 ;
      RECT 59.79 27.1 63.75 27.24 ;
      RECT 63.46 30.795 63.75 31.025 ;
      RECT 61.89 30.795 62.18 31.025 ;
      RECT 59.79 30.795 60.08 31.025 ;
      RECT 59.79 30.84 63.75 30.98 ;
      RECT 49.72 14.52 59.06 14.66 ;
      RECT 58.92 14.18 59.06 14.66 ;
      RECT 52.02 13.84 52.16 14.66 ;
      RECT 49.72 13.84 49.86 14.66 ;
      RECT 59.75 14.12 60.07 14.38 ;
      RECT 58.92 14.18 63.43 14.32 ;
      RECT 63.29 13.795 63.43 14.32 ;
      RECT 63.215 13.795 63.505 14.025 ;
      RECT 51.03 13.795 51.32 14.025 ;
      RECT 45.965 13.795 46.255 14.025 ;
      RECT 51.03 13.84 52.16 13.98 ;
      RECT 45.965 13.84 49.86 13.98 ;
      RECT 46.04 13.5 46.18 14.025 ;
      RECT 43.19 13.44 43.51 13.7 ;
      RECT 43.19 13.5 46.18 13.64 ;
      RECT 62.51 14.8 62.83 15.06 ;
      RECT 60.685 14.815 60.975 15.045 ;
      RECT 60.685 14.86 62.83 15 ;
      RECT 62.51 16.84 62.83 17.1 ;
      RECT 60.61 16.855 60.9 17.085 ;
      RECT 60.61 16.9 62.83 17.04 ;
      RECT 62.51 21.26 62.83 21.52 ;
      RECT 58.385 21.275 58.675 21.505 ;
      RECT 58.385 21.32 62.83 21.46 ;
      RECT 62.51 29.76 62.83 30.02 ;
      RECT 60.61 29.775 60.9 30.005 ;
      RECT 60.61 29.82 62.83 29.96 ;
      RECT 56.99 13.78 57.31 14.04 ;
      RECT 61.375 13.795 61.665 14.025 ;
      RECT 53.095 13.795 53.385 14.025 ;
      RECT 60.3 13.84 61.665 13.98 ;
      RECT 53.095 13.84 58.14 13.98 ;
      RECT 58 13.5 58.14 13.98 ;
      RECT 60.3 13.5 60.44 13.98 ;
      RECT 58 13.5 60.44 13.64 ;
      RECT 55.24 19.28 58.6 19.42 ;
      RECT 58.46 18.94 58.6 19.42 ;
      RECT 55.24 18.94 55.38 19.42 ;
      RECT 54.23 18.88 54.55 19.14 ;
      RECT 60.61 18.895 60.9 19.125 ;
      RECT 58.46 18.94 60.9 19.08 ;
      RECT 54.23 18.94 55.38 19.08 ;
      RECT 59.75 22.96 60.07 23.22 ;
      RECT 60.225 22.975 60.515 23.205 ;
      RECT 59.75 23.02 60.515 23.16 ;
      RECT 59.75 16.84 60.07 17.1 ;
      RECT 59.305 16.855 59.595 17.085 ;
      RECT 59.305 16.9 60.07 17.04 ;
      RECT 59.75 19.22 60.07 19.48 ;
      RECT 59.305 19.235 59.595 19.465 ;
      RECT 59.305 19.28 60.07 19.42 ;
      RECT 59.75 27.72 60.07 27.98 ;
      RECT 59.305 27.735 59.595 27.965 ;
      RECT 59.305 27.78 60.07 27.92 ;
      RECT 59.75 30.1 60.07 30.36 ;
      RECT 59.305 30.115 59.595 30.345 ;
      RECT 59.305 30.16 60.07 30.3 ;
      RECT 48.495 22.295 48.785 22.525 ;
      RECT 48.495 22.34 51.24 22.48 ;
      RECT 51.1 21.32 51.24 22.48 ;
      RECT 56.99 21.26 57.31 21.52 ;
      RECT 51.47 21.26 51.79 21.52 ;
      RECT 51.1 21.32 57.31 21.46 ;
      RECT 56.99 32.14 57.31 32.4 ;
      RECT 55.625 32.155 55.915 32.385 ;
      RECT 55.625 32.2 57.31 32.34 ;
      RECT 48.71 15.82 49.03 16.08 ;
      RECT 57.005 15.835 57.295 16.065 ;
      RECT 48.71 15.88 57.295 16.02 ;
      RECT 48.365 18.54 48.685 18.8 ;
      RECT 56.545 18.555 56.835 18.785 ;
      RECT 48.365 18.6 56.835 18.74 ;
      RECT 56.075 21.955 56.365 22.185 ;
      RECT 53.555 21.955 53.845 22.185 ;
      RECT 52.365 21.955 52.655 22.185 ;
      RECT 52.365 22 56.365 22.14 ;
      RECT 55.64 21.615 55.93 21.845 ;
      RECT 54.07 21.615 54.36 21.845 ;
      RECT 51.97 21.615 52.26 21.845 ;
      RECT 51.97 21.66 55.93 21.8 ;
      RECT 54.23 34.86 54.55 35.12 ;
      RECT 55.165 34.875 55.455 35.105 ;
      RECT 54.23 34.92 55.455 35.06 ;
      RECT 54.695 16.515 54.985 16.745 ;
      RECT 52.175 16.515 52.465 16.745 ;
      RECT 50.985 16.515 51.275 16.745 ;
      RECT 50.985 16.56 54.985 16.7 ;
      RECT 54.23 14.8 54.55 15.06 ;
      RECT 53.785 14.815 54.075 15.045 ;
      RECT 53.785 14.86 54.55 15 ;
      RECT 54.26 16.175 54.55 16.405 ;
      RECT 52.69 16.175 52.98 16.405 ;
      RECT 50.59 16.175 50.88 16.405 ;
      RECT 50.59 16.22 54.55 16.36 ;
      RECT 54.23 22.62 54.55 22.88 ;
      RECT 52.79 22.635 53.08 22.865 ;
      RECT 52.79 22.68 54.55 22.82 ;
      RECT 48.495 27.735 48.785 27.965 ;
      RECT 48.57 27.44 48.71 27.965 ;
      RECT 54.23 27.38 54.55 27.64 ;
      RECT 51.47 27.38 51.79 27.64 ;
      RECT 48.57 27.44 54.55 27.58 ;
      RECT 54.23 30.1 54.55 30.36 ;
      RECT 48.495 30.115 48.785 30.345 ;
      RECT 48.495 30.16 54.55 30.3 ;
      RECT 54.23 30.78 54.55 31.04 ;
      RECT 45.95 30.78 46.27 31.04 ;
      RECT 45.95 30.84 54.55 30.98 ;
      RECT 47.42 30.115 47.56 30.98 ;
      RECT 47.345 30.115 47.635 30.345 ;
      RECT 54.235 19.575 54.525 19.805 ;
      RECT 51.715 19.575 52.005 19.805 ;
      RECT 50.525 19.575 50.815 19.805 ;
      RECT 50.525 19.62 54.525 19.76 ;
      RECT 54.235 25.015 54.525 25.245 ;
      RECT 51.715 25.015 52.005 25.245 ;
      RECT 50.525 25.015 50.815 25.245 ;
      RECT 50.525 25.06 54.525 25.2 ;
      RECT 53.8 19.915 54.09 20.145 ;
      RECT 52.23 19.915 52.52 20.145 ;
      RECT 50.13 19.915 50.42 20.145 ;
      RECT 50.13 19.96 54.09 20.1 ;
      RECT 53.8 25.355 54.09 25.585 ;
      RECT 52.23 25.355 52.52 25.585 ;
      RECT 50.13 25.355 50.42 25.585 ;
      RECT 50.13 25.4 54.09 25.54 ;
      RECT 53.315 32.835 53.605 33.065 ;
      RECT 50.795 32.835 51.085 33.065 ;
      RECT 49.605 32.835 49.895 33.065 ;
      RECT 49.605 32.88 53.605 33.02 ;
      RECT 52.88 32.495 53.17 32.725 ;
      RECT 51.31 32.495 51.6 32.725 ;
      RECT 49.21 32.495 49.5 32.725 ;
      RECT 49.21 32.54 53.17 32.68 ;
      RECT 52.855 35.895 53.145 36.125 ;
      RECT 50.335 35.895 50.625 36.125 ;
      RECT 49.145 35.895 49.435 36.125 ;
      RECT 49.145 35.94 53.145 36.08 ;
      RECT 52.42 36.235 52.71 36.465 ;
      RECT 50.85 36.235 51.14 36.465 ;
      RECT 48.75 36.235 49.04 36.465 ;
      RECT 48.75 36.28 52.71 36.42 ;
      RECT 52.405 13.455 52.695 13.685 ;
      RECT 52.48 13.16 52.62 13.685 ;
      RECT 51.47 13.1 51.79 13.36 ;
      RECT 51.47 13.16 52.62 13.3 ;
      RECT 48.71 13.44 49.03 13.7 ;
      RECT 51.945 13.455 52.235 13.685 ;
      RECT 48.71 13.5 52.235 13.64 ;
      RECT 51.47 14.12 51.79 14.38 ;
      RECT 50.67 14.18 51.79 14.32 ;
      RECT 50.67 13.795 50.81 14.32 ;
      RECT 50.595 13.795 50.885 14.025 ;
      RECT 51.47 14.8 51.79 15.06 ;
      RECT 47.345 14.815 47.635 15.045 ;
      RECT 47.345 14.86 51.79 15 ;
      RECT 51.47 16.84 51.79 17.1 ;
      RECT 51.41 16.855 51.79 17.085 ;
      RECT 51.47 17.52 51.79 17.78 ;
      RECT 47.805 17.535 48.095 17.765 ;
      RECT 47.805 17.58 51.79 17.72 ;
      RECT 51.47 18.88 51.79 19.14 ;
      RECT 50.95 18.895 51.24 19.125 ;
      RECT 50.95 18.94 51.79 19.08 ;
      RECT 51.47 22.96 51.79 23.22 ;
      RECT 49.185 22.975 49.475 23.205 ;
      RECT 49.185 23.02 51.79 23.16 ;
      RECT 51.47 24.32 51.79 24.58 ;
      RECT 50.95 24.335 51.24 24.565 ;
      RECT 50.95 24.38 51.79 24.52 ;
      RECT 51.47 28.4 51.79 28.66 ;
      RECT 49.185 28.415 49.475 28.645 ;
      RECT 49.185 28.46 51.79 28.6 ;
      RECT 51.47 31.12 51.79 31.38 ;
      RECT 49.185 31.135 49.475 31.365 ;
      RECT 49.185 31.18 51.79 31.32 ;
      RECT 51.47 33.16 51.79 33.42 ;
      RECT 50.03 33.175 50.32 33.405 ;
      RECT 50.03 33.22 51.79 33.36 ;
      RECT 51.47 35.2 51.79 35.46 ;
      RECT 49.57 35.215 49.86 35.445 ;
      RECT 49.57 35.26 51.79 35.4 ;
      RECT 48.71 16.84 49.03 17.1 ;
      RECT 50.105 16.855 50.395 17.085 ;
      RECT 48.71 16.9 50.395 17.04 ;
      RECT 48.71 19.22 49.03 19.48 ;
      RECT 49.645 19.235 49.935 19.465 ;
      RECT 48.71 19.28 49.935 19.42 ;
      RECT 48.71 24.66 49.03 24.92 ;
      RECT 49.645 24.675 49.935 24.905 ;
      RECT 48.71 24.72 49.935 24.86 ;
      RECT 48.265 35.895 48.555 36.125 ;
      RECT 48.265 35.94 48.94 36.08 ;
      RECT 48.8 35.54 48.94 36.08 ;
      RECT 48.71 35.54 49.03 35.8 ;
      RECT 48.365 14.46 48.685 14.72 ;
      RECT 45.95 14.46 46.27 14.72 ;
      RECT 45.605 14.52 48.685 14.66 ;
      RECT 45.605 13.795 45.745 14.66 ;
      RECT 45.53 13.795 45.82 14.025 ;
      RECT 48.25 9.36 48.57 9.62 ;
      RECT 42.73 9.36 43.05 9.62 ;
      RECT 47.42 9.42 48.57 9.56 ;
      RECT 42.73 9.42 43.88 9.56 ;
      RECT 43.74 8.74 43.88 9.56 ;
      RECT 47.42 8.74 47.56 9.56 ;
      RECT 43.74 8.74 47.56 8.88 ;
      RECT 45.95 22.96 46.27 23.22 ;
      RECT 45.95 23.02 48.02 23.16 ;
      RECT 47.88 21.32 48.02 23.16 ;
      RECT 47.805 22.295 48.095 22.525 ;
      RECT 33.16 21.66 42.5 21.8 ;
      RECT 42.36 21.49 42.5 21.8 ;
      RECT 33.16 21.32 33.3 21.8 ;
      RECT 42.36 21.49 47.1 21.63 ;
      RECT 46.96 21.32 47.1 21.63 ;
      RECT 32.15 21.26 32.47 21.52 ;
      RECT 46.96 21.32 48.02 21.46 ;
      RECT 32.15 21.32 33.3 21.46 ;
      RECT 40.43 22.62 40.75 22.88 ;
      RECT 29.39 22.62 29.71 22.88 ;
      RECT 47.345 22.635 47.635 22.865 ;
      RECT 29.39 22.68 47.635 22.82 ;
      RECT 47.115 27.735 47.405 27.965 ;
      RECT 47.19 26.76 47.33 27.965 ;
      RECT 45.95 26.7 46.27 26.96 ;
      RECT 45.95 26.76 47.33 26.9 ;
      RECT 46.655 22.295 46.945 22.525 ;
      RECT 46.73 22 46.87 22.525 ;
      RECT 43.19 21.94 43.51 22.2 ;
      RECT 43.19 22 46.87 22.14 ;
      RECT 46.655 27.735 46.945 27.965 ;
      RECT 46.73 27.44 46.87 27.965 ;
      RECT 43.19 27.38 43.51 27.64 ;
      RECT 43.19 27.44 46.87 27.58 ;
      RECT 43.19 30.44 43.51 30.7 ;
      RECT 43.19 30.5 46.87 30.64 ;
      RECT 46.73 30.115 46.87 30.64 ;
      RECT 46.655 30.115 46.945 30.345 ;
      RECT 46.425 16.855 46.715 17.085 ;
      RECT 46.5 15.88 46.64 17.085 ;
      RECT 45.95 15.82 46.27 16.08 ;
      RECT 45.95 15.88 46.64 16.02 ;
      RECT 45.95 11.4 46.27 11.66 ;
      RECT 30.785 11.415 31.075 11.645 ;
      RECT 30.785 11.46 46.27 11.6 ;
      RECT 37.685 13.795 37.975 14.025 ;
      RECT 37.76 13.16 37.9 14.025 ;
      RECT 38.68 13.5 42.5 13.64 ;
      RECT 42.36 13.16 42.5 13.64 ;
      RECT 38.68 13.16 38.82 13.64 ;
      RECT 45.95 13.1 46.27 13.36 ;
      RECT 42.36 13.16 46.27 13.3 ;
      RECT 37.76 13.16 38.82 13.3 ;
      RECT 44.585 16.855 44.875 17.085 ;
      RECT 44.66 16.22 44.8 17.085 ;
      RECT 45.95 16.5 46.27 16.76 ;
      RECT 44.66 16.56 46.27 16.7 ;
      RECT 43.19 16.16 43.51 16.42 ;
      RECT 43.19 16.22 44.8 16.36 ;
      RECT 34.91 17.52 35.23 17.78 ;
      RECT 42.36 17.58 46.18 17.72 ;
      RECT 46.04 17.195 46.18 17.72 ;
      RECT 34.91 17.58 36.06 17.72 ;
      RECT 35.92 17.24 36.06 17.72 ;
      RECT 42.36 17.41 42.5 17.72 ;
      RECT 38.22 17.41 42.5 17.55 ;
      RECT 45.965 17.195 46.255 17.425 ;
      RECT 38.22 17.24 38.36 17.55 ;
      RECT 35.92 17.24 38.36 17.38 ;
      RECT 43.19 14.8 43.51 15.06 ;
      RECT 45.505 14.815 45.795 15.045 ;
      RECT 43.19 14.86 45.795 15 ;
      RECT 43.19 17.18 43.51 17.44 ;
      RECT 43.19 17.24 45.49 17.38 ;
      RECT 45.35 16.855 45.49 17.38 ;
      RECT 45.275 16.855 45.565 17.085 ;
      RECT 34.91 14.8 35.23 15.06 ;
      RECT 34.91 14.86 35.6 15 ;
      RECT 35.46 13.84 35.6 15 ;
      RECT 43.19 14.12 43.51 14.38 ;
      RECT 35.46 14.18 43.51 14.32 ;
      RECT 20.205 13.795 20.495 14.025 ;
      RECT 20.205 13.84 35.6 13.98 ;
      RECT 32.15 17.18 32.47 17.44 ;
      RECT 30.86 17.24 32.47 17.38 ;
      RECT 30.86 16.855 31 17.38 ;
      RECT 30.785 16.855 31.075 17.085 ;
      RECT 29.39 17.18 29.71 17.44 ;
      RECT 28.56 17.24 29.71 17.38 ;
      RECT 20.28 17.24 22.26 17.38 ;
      RECT 22.12 16.9 22.26 17.38 ;
      RECT 28.56 16.9 28.7 17.38 ;
      RECT 20.28 16.855 20.42 17.38 ;
      RECT 20.205 16.855 20.495 17.085 ;
      RECT 22.12 16.9 28.7 17.04 ;
      RECT 183.95 21.26 184.27 21.52 ;
      RECT 181.19 24.66 181.51 24.92 ;
      RECT 172.91 22.62 173.23 22.88 ;
      RECT 153.59 16.84 153.91 17.1 ;
      RECT 153.59 21.94 153.91 22.2 ;
      RECT 142.55 16.84 142.87 17.1 ;
      RECT 98.39 11.4 98.71 11.66 ;
      RECT 95.63 30.1 95.95 30.36 ;
      RECT 62.51 11.4 62.83 11.66 ;
      RECT 62.51 13.78 62.83 14.04 ;
      RECT 48.71 32.82 49.03 33.08 ;
      RECT 45.95 22.28 46.27 22.54 ;
      RECT 45.95 27.72 46.27 27.98 ;
      RECT 45.95 30.1 46.27 30.36 ;
      RECT 40.43 16.84 40.75 17.1 ;
    LAYER via ;
      RECT 184.035 13.495 184.185 13.645 ;
      RECT 184.035 21.315 184.185 21.465 ;
      RECT 181.275 24.715 181.425 24.865 ;
      RECT 181.275 28.115 181.425 28.265 ;
      RECT 175.755 14.515 175.905 14.665 ;
      RECT 175.755 15.875 175.905 16.025 ;
      RECT 175.755 16.895 175.905 17.045 ;
      RECT 175.755 21.315 175.905 21.465 ;
      RECT 175.755 22.675 175.905 22.825 ;
      RECT 175.755 24.035 175.905 24.185 ;
      RECT 172.995 10.435 173.145 10.585 ;
      RECT 172.995 19.955 173.145 20.105 ;
      RECT 172.995 22.675 173.145 22.825 ;
      RECT 172.995 24.035 173.145 24.185 ;
      RECT 172.995 24.715 173.145 24.865 ;
      RECT 170.235 17.235 170.385 17.385 ;
      RECT 170.235 21.655 170.385 21.805 ;
      RECT 167.475 12.135 167.625 12.285 ;
      RECT 167.475 13.495 167.625 13.645 ;
      RECT 167.475 14.855 167.625 15.005 ;
      RECT 167.475 18.595 167.625 18.745 ;
      RECT 167.475 20.295 167.625 20.445 ;
      RECT 167.475 24.375 167.625 24.525 ;
      RECT 167.475 25.395 167.625 25.545 ;
      RECT 167.475 26.755 167.625 26.905 ;
      RECT 164.715 19.275 164.865 19.425 ;
      RECT 164.715 23.015 164.865 23.165 ;
      RECT 164.715 24.035 164.865 24.185 ;
      RECT 161.955 22.335 162.105 22.485 ;
      RECT 161.955 23.015 162.105 23.165 ;
      RECT 161.955 26.755 162.105 26.905 ;
      RECT 159.195 13.835 159.345 13.985 ;
      RECT 159.195 22.335 159.345 22.485 ;
      RECT 159.195 27.775 159.345 27.925 ;
      RECT 156.435 16.895 156.585 17.045 ;
      RECT 156.435 23.015 156.585 23.165 ;
      RECT 156.435 28.115 156.585 28.265 ;
      RECT 156.435 30.155 156.585 30.305 ;
      RECT 153.675 16.895 153.825 17.045 ;
      RECT 153.675 19.275 153.825 19.425 ;
      RECT 153.675 21.995 153.825 22.145 ;
      RECT 153.675 22.675 153.825 22.825 ;
      RECT 153.675 24.035 153.825 24.185 ;
      RECT 153.675 25.395 153.825 25.545 ;
      RECT 153.675 26.755 153.825 26.905 ;
      RECT 150.915 16.555 151.065 16.705 ;
      RECT 150.915 25.735 151.065 25.885 ;
      RECT 150.915 27.775 151.065 27.925 ;
      RECT 150.915 29.815 151.065 29.965 ;
      RECT 148.155 11.455 148.305 11.605 ;
      RECT 148.155 16.895 148.305 17.045 ;
      RECT 148.155 17.575 148.305 17.725 ;
      RECT 148.155 18.935 148.305 19.085 ;
      RECT 148.155 19.615 148.305 19.765 ;
      RECT 148.155 22.335 148.305 22.485 ;
      RECT 148.155 24.035 148.305 24.185 ;
      RECT 145.395 13.835 145.545 13.985 ;
      RECT 145.395 16.215 145.545 16.365 ;
      RECT 145.395 17.575 145.545 17.725 ;
      RECT 145.395 18.595 145.545 18.745 ;
      RECT 145.395 24.375 145.545 24.525 ;
      RECT 145.395 26.755 145.545 26.905 ;
      RECT 142.635 16.215 142.785 16.365 ;
      RECT 142.635 16.895 142.785 17.045 ;
      RECT 142.635 17.575 142.785 17.725 ;
      RECT 142.635 18.595 142.785 18.745 ;
      RECT 142.635 19.275 142.785 19.425 ;
      RECT 142.635 19.955 142.785 20.105 ;
      RECT 142.635 24.715 142.785 24.865 ;
      RECT 142.635 25.395 142.785 25.545 ;
      RECT 142.635 27.095 142.785 27.245 ;
      RECT 142.635 29.475 142.785 29.625 ;
      RECT 142.635 31.175 142.785 31.325 ;
      RECT 139.875 11.455 140.025 11.605 ;
      RECT 139.875 17.575 140.025 17.725 ;
      RECT 139.875 23.015 140.025 23.165 ;
      RECT 139.875 29.815 140.025 29.965 ;
      RECT 137.115 13.495 137.265 13.645 ;
      RECT 137.115 17.575 137.265 17.725 ;
      RECT 137.115 18.595 137.265 18.745 ;
      RECT 137.115 22.675 137.265 22.825 ;
      RECT 137.115 24.035 137.265 24.185 ;
      RECT 137.115 24.715 137.265 24.865 ;
      RECT 137.115 28.115 137.265 28.265 ;
      RECT 137.115 29.475 137.265 29.625 ;
      RECT 137.115 30.155 137.265 30.305 ;
      RECT 134.355 14.855 134.505 15.005 ;
      RECT 134.355 16.555 134.505 16.705 ;
      RECT 134.355 20.295 134.505 20.445 ;
      RECT 134.355 23.015 134.505 23.165 ;
      RECT 134.355 27.435 134.505 27.585 ;
      RECT 131.595 14.175 131.745 14.325 ;
      RECT 131.595 16.895 131.745 17.045 ;
      RECT 131.595 17.575 131.745 17.725 ;
      RECT 131.595 18.935 131.745 19.085 ;
      RECT 131.595 21.315 131.745 21.465 ;
      RECT 131.595 25.055 131.745 25.205 ;
      RECT 131.595 27.775 131.745 27.925 ;
      RECT 128.835 13.835 128.985 13.985 ;
      RECT 128.835 14.515 128.985 14.665 ;
      RECT 128.835 16.215 128.985 16.365 ;
      RECT 128.835 16.895 128.985 17.045 ;
      RECT 128.835 18.595 128.985 18.745 ;
      RECT 128.835 19.275 128.985 19.425 ;
      RECT 128.835 19.955 128.985 20.105 ;
      RECT 128.835 22.335 128.985 22.485 ;
      RECT 128.835 24.035 128.985 24.185 ;
      RECT 126.075 11.455 126.225 11.605 ;
      RECT 126.075 16.215 126.225 16.365 ;
      RECT 126.075 16.895 126.225 17.045 ;
      RECT 126.075 17.575 126.225 17.725 ;
      RECT 126.075 21.315 126.225 21.465 ;
      RECT 126.075 22.675 126.225 22.825 ;
      RECT 126.075 24.715 126.225 24.865 ;
      RECT 126.075 26.755 126.225 26.905 ;
      RECT 126.075 29.475 126.225 29.625 ;
      RECT 126.075 30.495 126.225 30.645 ;
      RECT 123.315 12.135 123.465 12.285 ;
      RECT 123.315 13.495 123.465 13.645 ;
      RECT 123.315 14.855 123.465 15.005 ;
      RECT 123.315 16.215 123.465 16.365 ;
      RECT 123.315 17.235 123.465 17.385 ;
      RECT 123.315 18.595 123.465 18.745 ;
      RECT 123.315 19.275 123.465 19.425 ;
      RECT 123.315 22.335 123.465 22.485 ;
      RECT 123.315 27.435 123.465 27.585 ;
      RECT 123.315 28.115 123.465 28.265 ;
      RECT 123.315 30.155 123.465 30.305 ;
      RECT 123.315 32.195 123.465 32.345 ;
      RECT 120.555 13.155 120.705 13.305 ;
      RECT 120.555 18.935 120.705 19.085 ;
      RECT 120.555 27.095 120.705 27.245 ;
      RECT 120.555 27.775 120.705 27.925 ;
      RECT 120.555 30.155 120.705 30.305 ;
      RECT 118.195 14.515 118.345 14.665 ;
      RECT 118.195 16.215 118.345 16.365 ;
      RECT 117.795 12.135 117.945 12.285 ;
      RECT 117.795 13.835 117.945 13.985 ;
      RECT 117.795 16.895 117.945 17.045 ;
      RECT 117.795 18.935 117.945 19.085 ;
      RECT 117.795 19.615 117.945 19.765 ;
      RECT 117.795 22.335 117.945 22.485 ;
      RECT 117.795 24.715 117.945 24.865 ;
      RECT 117.795 25.735 117.945 25.885 ;
      RECT 117.795 28.115 117.945 28.265 ;
      RECT 117.795 38.315 117.945 38.465 ;
      RECT 115.035 18.595 115.185 18.745 ;
      RECT 115.035 19.275 115.185 19.425 ;
      RECT 115.035 21.315 115.185 21.465 ;
      RECT 115.035 29.475 115.185 29.625 ;
      RECT 112.275 13.835 112.425 13.985 ;
      RECT 112.275 15.875 112.425 16.025 ;
      RECT 112.275 16.895 112.425 17.045 ;
      RECT 112.275 17.575 112.425 17.725 ;
      RECT 112.275 22.675 112.425 22.825 ;
      RECT 112.275 24.035 112.425 24.185 ;
      RECT 112.275 25.735 112.425 25.885 ;
      RECT 112.275 27.095 112.425 27.245 ;
      RECT 112.275 27.775 112.425 27.925 ;
      RECT 112.275 30.155 112.425 30.305 ;
      RECT 112.275 30.835 112.425 30.985 ;
      RECT 112.275 32.195 112.425 32.345 ;
      RECT 109.515 14.515 109.665 14.665 ;
      RECT 109.515 15.875 109.665 16.025 ;
      RECT 109.515 17.575 109.665 17.725 ;
      RECT 109.515 24.715 109.665 24.865 ;
      RECT 109.515 27.775 109.665 27.925 ;
      RECT 109.515 29.475 109.665 29.625 ;
      RECT 103.995 15.875 104.145 16.025 ;
      RECT 103.995 17.575 104.145 17.725 ;
      RECT 101.235 16.895 101.385 17.045 ;
      RECT 101.235 21.315 101.385 21.465 ;
      RECT 101.235 22.675 101.385 22.825 ;
      RECT 101.235 29.475 101.385 29.625 ;
      RECT 98.475 11.455 98.625 11.605 ;
      RECT 98.475 13.155 98.625 13.305 ;
      RECT 98.475 24.035 98.625 24.185 ;
      RECT 98.475 28.115 98.625 28.265 ;
      RECT 95.715 13.155 95.865 13.305 ;
      RECT 95.715 13.835 95.865 13.985 ;
      RECT 95.715 16.895 95.865 17.045 ;
      RECT 95.715 18.935 95.865 19.085 ;
      RECT 95.715 20.295 95.865 20.445 ;
      RECT 95.715 24.035 95.865 24.185 ;
      RECT 95.715 29.475 95.865 29.625 ;
      RECT 95.715 30.155 95.865 30.305 ;
      RECT 92.955 13.155 93.105 13.305 ;
      RECT 92.955 16.555 93.105 16.705 ;
      RECT 92.955 17.575 93.105 17.725 ;
      RECT 92.955 18.935 93.105 19.085 ;
      RECT 92.955 19.615 93.105 19.765 ;
      RECT 92.955 22.335 93.105 22.485 ;
      RECT 92.955 23.015 93.105 23.165 ;
      RECT 92.955 27.095 93.105 27.245 ;
      RECT 92.955 27.775 93.105 27.925 ;
      RECT 92.955 29.815 93.105 29.965 ;
      RECT 90.195 11.455 90.345 11.605 ;
      RECT 90.195 14.515 90.345 14.665 ;
      RECT 90.195 18.935 90.345 19.085 ;
      RECT 90.195 21.315 90.345 21.465 ;
      RECT 90.195 22.335 90.345 22.485 ;
      RECT 90.195 24.715 90.345 24.865 ;
      RECT 90.195 28.455 90.345 28.605 ;
      RECT 90.195 29.815 90.345 29.965 ;
      RECT 87.435 11.795 87.585 11.945 ;
      RECT 87.435 14.855 87.585 15.005 ;
      RECT 87.435 15.875 87.585 16.025 ;
      RECT 87.435 16.895 87.585 17.045 ;
      RECT 87.435 18.595 87.585 18.745 ;
      RECT 87.435 19.615 87.585 19.765 ;
      RECT 87.435 31.175 87.585 31.325 ;
      RECT 84.675 16.215 84.825 16.365 ;
      RECT 84.675 18.595 84.825 18.745 ;
      RECT 84.675 20.295 84.825 20.445 ;
      RECT 84.675 21.315 84.825 21.465 ;
      RECT 84.675 24.035 84.825 24.185 ;
      RECT 84.675 27.435 84.825 27.585 ;
      RECT 84.675 29.475 84.825 29.625 ;
      RECT 84.675 30.495 84.825 30.645 ;
      RECT 84.675 32.195 84.825 32.345 ;
      RECT 82.3 13.835 82.45 13.985 ;
      RECT 81.915 11.455 82.065 11.605 ;
      RECT 81.915 16.215 82.065 16.365 ;
      RECT 81.915 17.575 82.065 17.725 ;
      RECT 81.915 18.935 82.065 19.085 ;
      RECT 81.915 19.615 82.065 19.765 ;
      RECT 81.915 23.015 82.065 23.165 ;
      RECT 81.915 30.835 82.065 30.985 ;
      RECT 81.915 32.195 82.065 32.345 ;
      RECT 79.155 16.895 79.305 17.045 ;
      RECT 79.155 17.575 79.305 17.725 ;
      RECT 79.155 18.935 79.305 19.085 ;
      RECT 79.155 20.295 79.305 20.445 ;
      RECT 79.155 24.375 79.305 24.525 ;
      RECT 79.155 29.475 79.305 29.625 ;
      RECT 79.155 30.155 79.305 30.305 ;
      RECT 76.395 23.015 76.545 23.165 ;
      RECT 76.395 29.475 76.545 29.625 ;
      RECT 76.395 30.155 76.545 30.305 ;
      RECT 76.395 31.175 76.545 31.325 ;
      RECT 76.395 32.535 76.545 32.685 ;
      RECT 73.635 11.455 73.785 11.605 ;
      RECT 73.635 13.155 73.785 13.305 ;
      RECT 73.635 15.875 73.785 16.025 ;
      RECT 73.635 16.555 73.785 16.705 ;
      RECT 73.635 17.575 73.785 17.725 ;
      RECT 73.635 18.595 73.785 18.745 ;
      RECT 73.635 19.275 73.785 19.425 ;
      RECT 73.635 25.055 73.785 25.205 ;
      RECT 73.635 27.095 73.785 27.245 ;
      RECT 73.635 27.775 73.785 27.925 ;
      RECT 73.635 28.455 73.785 28.605 ;
      RECT 73.635 29.475 73.785 29.625 ;
      RECT 73.635 30.155 73.785 30.305 ;
      RECT 73.635 30.835 73.785 30.985 ;
      RECT 73.635 32.195 73.785 32.345 ;
      RECT 70.875 13.835 71.025 13.985 ;
      RECT 70.875 16.215 71.025 16.365 ;
      RECT 70.875 17.575 71.025 17.725 ;
      RECT 70.875 31.175 71.025 31.325 ;
      RECT 68.115 14.855 68.265 15.005 ;
      RECT 68.115 16.555 68.265 16.705 ;
      RECT 68.115 17.575 68.265 17.725 ;
      RECT 68.115 24.035 68.265 24.185 ;
      RECT 68.115 27.775 68.265 27.925 ;
      RECT 65.355 12.135 65.505 12.285 ;
      RECT 65.355 15.875 65.505 16.025 ;
      RECT 65.355 19.615 65.505 19.765 ;
      RECT 65.355 22.335 65.505 22.485 ;
      RECT 65.355 27.435 65.505 27.585 ;
      RECT 65.355 32.535 65.505 32.685 ;
      RECT 62.595 11.455 62.745 11.605 ;
      RECT 62.595 13.155 62.745 13.305 ;
      RECT 62.595 13.835 62.745 13.985 ;
      RECT 62.595 14.855 62.745 15.005 ;
      RECT 62.595 16.895 62.745 17.045 ;
      RECT 62.595 18.595 62.745 18.745 ;
      RECT 62.595 21.315 62.745 21.465 ;
      RECT 62.595 25.395 62.745 25.545 ;
      RECT 62.595 26.755 62.745 26.905 ;
      RECT 62.595 28.455 62.745 28.605 ;
      RECT 62.595 29.815 62.745 29.965 ;
      RECT 59.835 14.175 59.985 14.325 ;
      RECT 59.835 16.895 59.985 17.045 ;
      RECT 59.835 19.275 59.985 19.425 ;
      RECT 59.835 23.015 59.985 23.165 ;
      RECT 59.835 27.775 59.985 27.925 ;
      RECT 59.835 30.155 59.985 30.305 ;
      RECT 57.075 13.835 57.225 13.985 ;
      RECT 57.075 17.235 57.225 17.385 ;
      RECT 57.075 18.595 57.225 18.745 ;
      RECT 57.075 21.315 57.225 21.465 ;
      RECT 57.075 28.115 57.225 28.265 ;
      RECT 57.075 32.195 57.225 32.345 ;
      RECT 54.315 14.855 54.465 15.005 ;
      RECT 54.315 18.935 54.465 19.085 ;
      RECT 54.315 20.295 54.465 20.445 ;
      RECT 54.315 22.675 54.465 22.825 ;
      RECT 54.315 27.435 54.465 27.585 ;
      RECT 54.315 30.155 54.465 30.305 ;
      RECT 54.315 30.835 54.465 30.985 ;
      RECT 54.315 34.915 54.465 35.065 ;
      RECT 51.555 12.135 51.705 12.285 ;
      RECT 51.555 13.155 51.705 13.305 ;
      RECT 51.555 14.175 51.705 14.325 ;
      RECT 51.555 14.855 51.705 15.005 ;
      RECT 51.555 16.895 51.705 17.045 ;
      RECT 51.555 17.575 51.705 17.725 ;
      RECT 51.555 18.935 51.705 19.085 ;
      RECT 51.555 21.315 51.705 21.465 ;
      RECT 51.555 23.015 51.705 23.165 ;
      RECT 51.555 24.375 51.705 24.525 ;
      RECT 51.555 27.435 51.705 27.585 ;
      RECT 51.555 28.455 51.705 28.605 ;
      RECT 51.555 31.175 51.705 31.325 ;
      RECT 51.555 33.215 51.705 33.365 ;
      RECT 51.555 35.255 51.705 35.405 ;
      RECT 48.795 13.495 48.945 13.645 ;
      RECT 48.795 15.875 48.945 16.025 ;
      RECT 48.795 16.895 48.945 17.045 ;
      RECT 48.795 19.275 48.945 19.425 ;
      RECT 48.795 24.715 48.945 24.865 ;
      RECT 48.795 32.875 48.945 33.025 ;
      RECT 48.795 35.595 48.945 35.745 ;
      RECT 48.45 14.515 48.6 14.665 ;
      RECT 48.45 18.595 48.6 18.745 ;
      RECT 48.335 9.415 48.485 9.565 ;
      RECT 46.035 11.455 46.185 11.605 ;
      RECT 46.035 13.155 46.185 13.305 ;
      RECT 46.035 14.515 46.185 14.665 ;
      RECT 46.035 15.875 46.185 16.025 ;
      RECT 46.035 16.555 46.185 16.705 ;
      RECT 46.035 22.335 46.185 22.485 ;
      RECT 46.035 23.015 46.185 23.165 ;
      RECT 46.035 24.375 46.185 24.525 ;
      RECT 46.035 26.755 46.185 26.905 ;
      RECT 46.035 27.775 46.185 27.925 ;
      RECT 46.035 29.475 46.185 29.625 ;
      RECT 46.035 30.155 46.185 30.305 ;
      RECT 46.035 30.835 46.185 30.985 ;
      RECT 43.275 13.495 43.425 13.645 ;
      RECT 43.275 14.175 43.425 14.325 ;
      RECT 43.275 14.855 43.425 15.005 ;
      RECT 43.275 16.215 43.425 16.365 ;
      RECT 43.275 17.235 43.425 17.385 ;
      RECT 43.275 21.995 43.425 22.145 ;
      RECT 43.275 27.435 43.425 27.585 ;
      RECT 43.275 30.495 43.425 30.645 ;
      RECT 42.815 9.415 42.965 9.565 ;
      RECT 40.515 16.895 40.665 17.045 ;
      RECT 40.515 22.675 40.665 22.825 ;
      RECT 40.515 29.815 40.665 29.965 ;
      RECT 40.515 38.315 40.665 38.465 ;
      RECT 34.995 14.855 35.145 15.005 ;
      RECT 34.995 17.575 35.145 17.725 ;
      RECT 32.235 17.235 32.385 17.385 ;
      RECT 32.235 21.315 32.385 21.465 ;
      RECT 29.475 17.235 29.625 17.385 ;
      RECT 29.475 22.675 29.625 22.825 ;
    LAYER met2 ;
      RECT 183.98 21.23 184.24 21.55 ;
      RECT 184.04 13.41 184.18 21.55 ;
      RECT 183.98 13.41 184.24 13.73 ;
      RECT 181.22 28.03 181.48 28.35 ;
      RECT 181.28 24.63 181.42 28.35 ;
      RECT 181.22 24.63 181.48 24.95 ;
      RECT 175.7 15.79 175.96 16.11 ;
      RECT 175.76 14.43 175.9 16.11 ;
      RECT 175.7 14.43 175.96 14.75 ;
      RECT 175.7 21.23 175.96 21.55 ;
      RECT 175.76 16.81 175.9 21.55 ;
      RECT 175.7 16.81 175.96 17.13 ;
      RECT 175.7 23.95 175.96 24.27 ;
      RECT 175.76 22.59 175.9 24.27 ;
      RECT 175.7 22.59 175.96 22.91 ;
      RECT 172.94 24.63 173.2 24.95 ;
      RECT 172.94 24.72 173.6 24.86 ;
      RECT 173.46 22.68 173.6 24.86 ;
      RECT 172.94 22.59 173.2 22.91 ;
      RECT 172.94 22.68 173.6 22.82 ;
      RECT 172.94 23.95 173.2 24.27 ;
      RECT 172.54 24.04 173.2 24.18 ;
      RECT 172.54 22 172.68 24.18 ;
      RECT 172.54 22 173.14 22.14 ;
      RECT 173 19.87 173.14 22.14 ;
      RECT 172.94 19.87 173.2 20.19 ;
      RECT 172.54 19.96 173.2 20.1 ;
      RECT 172.54 18.26 172.68 20.1 ;
      RECT 172.54 18.26 172.91 18.4 ;
      RECT 172.77 14.86 172.91 18.4 ;
      RECT 172.54 14.86 172.91 15 ;
      RECT 172.54 10.44 172.68 15 ;
      RECT 172.94 10.35 173.2 10.67 ;
      RECT 172.54 10.44 173.2 10.58 ;
      RECT 170.18 21.57 170.44 21.89 ;
      RECT 170.24 17.15 170.38 21.89 ;
      RECT 170.17 18.525 170.45 18.895 ;
      RECT 170.18 17.15 170.44 17.47 ;
      RECT 167.42 13.41 167.68 13.73 ;
      RECT 167.48 12.05 167.62 13.73 ;
      RECT 167.42 12.05 167.68 12.37 ;
      RECT 167.42 18.51 167.68 18.83 ;
      RECT 167.48 14.77 167.62 18.83 ;
      RECT 167.42 14.77 167.68 15.09 ;
      RECT 167.42 24.29 167.68 24.61 ;
      RECT 167.48 20.21 167.62 24.61 ;
      RECT 167.42 20.21 167.68 20.53 ;
      RECT 167.42 26.67 167.68 26.99 ;
      RECT 167.48 25.31 167.62 26.99 ;
      RECT 167.42 25.31 167.68 25.63 ;
      RECT 164.66 19.19 164.92 19.51 ;
      RECT 164.72 18.525 164.86 19.51 ;
      RECT 164.65 18.525 164.93 18.895 ;
      RECT 164.65 25.845 164.93 26.215 ;
      RECT 164.72 22.93 164.86 26.215 ;
      RECT 164.66 23.95 164.92 24.27 ;
      RECT 164.66 22.93 164.92 23.25 ;
      RECT 161.9 22.25 162.16 22.57 ;
      RECT 161.96 18.525 162.1 22.57 ;
      RECT 161.89 18.525 162.17 18.895 ;
      RECT 161.9 26.67 162.16 26.99 ;
      RECT 161.96 22.93 162.1 26.99 ;
      RECT 161.9 22.93 162.16 23.25 ;
      RECT 159.14 27.69 159.4 28.01 ;
      RECT 159.2 13.75 159.34 28.01 ;
      RECT 159.14 22.25 159.4 22.57 ;
      RECT 159.14 13.75 159.4 14.07 ;
      RECT 156.38 30.07 156.64 30.39 ;
      RECT 156.44 16.81 156.58 30.39 ;
      RECT 156.38 28.03 156.64 28.35 ;
      RECT 156.38 22.93 156.64 23.25 ;
      RECT 156.38 16.81 156.64 17.13 ;
      RECT 153.62 21.91 153.88 22.23 ;
      RECT 153.68 16.81 153.82 22.23 ;
      RECT 153.62 19.19 153.88 19.51 ;
      RECT 153.61 18.525 153.89 18.895 ;
      RECT 153.62 16.81 153.88 17.13 ;
      RECT 153.62 23.95 153.88 24.27 ;
      RECT 153.68 22.59 153.82 24.27 ;
      RECT 153.62 22.59 153.88 22.91 ;
      RECT 153.62 26.67 153.88 26.99 ;
      RECT 153.68 25.31 153.82 26.99 ;
      RECT 153.62 25.31 153.88 25.63 ;
      RECT 150.86 16.47 151.12 16.79 ;
      RECT 150.46 16.56 151.12 16.7 ;
      RECT 150.46 15.54 150.6 16.7 ;
      RECT 150.46 15.54 150.83 15.68 ;
      RECT 150.69 10.44 150.83 15.68 ;
      RECT 150.46 10.44 150.83 10.58 ;
      RECT 150.46 9.375 150.6 10.58 ;
      RECT 150.39 9.375 150.67 9.745 ;
      RECT 150.86 29.73 151.12 30.05 ;
      RECT 150.92 25.65 151.06 30.05 ;
      RECT 150.86 27.69 151.12 28.01 ;
      RECT 150.86 25.65 151.12 25.97 ;
      RECT 148.1 23.95 148.36 24.27 ;
      RECT 148.16 21.32 148.3 24.27 ;
      RECT 148.1 22.25 148.36 22.57 ;
      RECT 148.16 21.32 148.76 21.46 ;
      RECT 148.62 16.9 148.76 21.46 ;
      RECT 148.07 16.84 148.39 17.1 ;
      RECT 148.07 16.9 148.76 17.04 ;
      RECT 148.1 19.53 148.36 19.85 ;
      RECT 147.7 19.62 148.36 19.76 ;
      RECT 147.7 16.56 147.84 19.76 ;
      RECT 147.7 16.56 148.3 16.7 ;
      RECT 148.16 11.37 148.3 16.7 ;
      RECT 148.1 11.37 148.36 11.69 ;
      RECT 148.1 18.85 148.36 19.17 ;
      RECT 148.16 17.49 148.3 19.17 ;
      RECT 148.1 17.49 148.36 17.81 ;
      RECT 145.34 16.13 145.6 16.45 ;
      RECT 145.4 13.75 145.54 16.45 ;
      RECT 145.34 13.75 145.6 14.07 ;
      RECT 145.34 18.51 145.6 18.83 ;
      RECT 145.4 17.49 145.54 18.83 ;
      RECT 145.34 17.49 145.6 17.81 ;
      RECT 145.34 26.67 145.6 26.99 ;
      RECT 145.4 24.29 145.54 26.99 ;
      RECT 145.34 24.29 145.6 24.61 ;
      RECT 142.58 31.09 142.84 31.41 ;
      RECT 142.64 25.31 142.78 31.41 ;
      RECT 142.58 29.39 142.84 29.71 ;
      RECT 142.58 27.01 142.84 27.33 ;
      RECT 142.58 25.31 142.84 25.63 ;
      RECT 142.58 25.4 143.24 25.54 ;
      RECT 143.1 14.98 143.24 25.54 ;
      RECT 142.58 19.87 142.84 20.19 ;
      RECT 142.58 19.96 143.24 20.1 ;
      RECT 142.58 16.13 142.84 16.45 ;
      RECT 142.64 14.865 142.78 16.45 ;
      RECT 142.57 14.865 142.85 15.235 ;
      RECT 142.57 14.98 143.24 15.12 ;
      RECT 142.57 18.525 142.85 18.895 ;
      RECT 142.58 18.51 142.84 18.895 ;
      RECT 142.64 17.49 142.78 18.895 ;
      RECT 142.58 17.49 142.84 17.81 ;
      RECT 142.58 24.63 142.84 24.95 ;
      RECT 142.18 24.72 142.84 24.86 ;
      RECT 142.18 16.9 142.32 24.86 ;
      RECT 142.58 19.19 142.84 19.51 ;
      RECT 142.18 19.28 142.84 19.42 ;
      RECT 142.58 16.81 142.84 17.13 ;
      RECT 142.18 16.9 142.84 17.04 ;
      RECT 139.82 17.49 140.08 17.81 ;
      RECT 139.82 17.58 140.48 17.72 ;
      RECT 140.34 9.375 140.48 17.72 ;
      RECT 140.27 9.375 140.55 9.745 ;
      RECT 139.82 29.73 140.08 30.05 ;
      RECT 139.88 18.6 140.02 30.05 ;
      RECT 139.82 22.93 140.08 23.25 ;
      RECT 139.42 18.6 140.02 18.74 ;
      RECT 139.42 16.56 139.56 18.74 ;
      RECT 139.42 16.56 139.79 16.7 ;
      RECT 139.65 12.48 139.79 16.7 ;
      RECT 139.65 12.48 140.02 12.62 ;
      RECT 139.88 11.37 140.02 12.62 ;
      RECT 139.82 11.37 140.08 11.69 ;
      RECT 137.06 18.51 137.32 18.83 ;
      RECT 137.12 13.41 137.26 18.83 ;
      RECT 137.06 17.49 137.32 17.81 ;
      RECT 137.06 13.41 137.32 13.73 ;
      RECT 137.06 23.95 137.32 24.27 ;
      RECT 137.12 22.59 137.26 24.27 ;
      RECT 137.06 22.59 137.32 22.91 ;
      RECT 137.06 30.07 137.32 30.39 ;
      RECT 136.66 30.16 137.32 30.3 ;
      RECT 136.66 27.44 136.8 30.3 ;
      RECT 136.66 27.44 137.26 27.58 ;
      RECT 137.12 24.63 137.26 27.58 ;
      RECT 137.06 24.63 137.32 24.95 ;
      RECT 137.06 29.39 137.32 29.71 ;
      RECT 137.12 28.03 137.26 29.71 ;
      RECT 137.06 28.03 137.32 28.35 ;
      RECT 134.3 20.21 134.56 20.53 ;
      RECT 134.36 14.77 134.5 20.53 ;
      RECT 134.3 16.47 134.56 16.79 ;
      RECT 134.3 14.77 134.56 15.09 ;
      RECT 134.3 27.35 134.56 27.67 ;
      RECT 134.36 22.93 134.5 27.67 ;
      RECT 134.3 22.93 134.56 23.25 ;
      RECT 131.54 24.97 131.8 25.29 ;
      RECT 131.6 23.36 131.74 25.29 ;
      RECT 131.6 23.36 132.2 23.5 ;
      RECT 132.06 21.32 132.2 23.5 ;
      RECT 131.54 21.23 131.8 21.55 ;
      RECT 131.54 21.32 132.2 21.46 ;
      RECT 131.54 16.81 131.8 17.13 ;
      RECT 131.6 14.09 131.74 17.13 ;
      RECT 131.53 14.865 131.81 15.235 ;
      RECT 131.54 14.09 131.8 14.41 ;
      RECT 131.54 27.69 131.8 28.01 ;
      RECT 131.6 25.845 131.74 28.01 ;
      RECT 131.53 25.845 131.81 26.215 ;
      RECT 131.54 18.85 131.8 19.17 ;
      RECT 131.6 17.49 131.74 19.17 ;
      RECT 131.54 17.49 131.8 17.81 ;
      RECT 128.78 18.51 129.04 18.83 ;
      RECT 128.78 18.6 129.44 18.74 ;
      RECT 129.3 14.52 129.44 18.74 ;
      RECT 128.75 16.16 129.07 16.42 ;
      RECT 128.84 15.88 128.98 16.42 ;
      RECT 128.84 15.88 129.44 16.02 ;
      RECT 128.78 14.43 129.04 14.75 ;
      RECT 128.78 14.52 129.44 14.66 ;
      RECT 128.78 23.95 129.04 24.27 ;
      RECT 128.38 24.04 129.04 24.18 ;
      RECT 128.38 13.84 128.52 24.18 ;
      RECT 128.78 19.19 129.04 19.51 ;
      RECT 128.38 19.28 129.04 19.42 ;
      RECT 128.77 17.915 129.05 18.285 ;
      RECT 128.38 17.92 129.05 18.06 ;
      RECT 128.84 16.81 128.98 18.285 ;
      RECT 128.78 16.81 129.04 17.13 ;
      RECT 128.78 13.75 129.04 14.07 ;
      RECT 128.38 13.84 129.04 13.98 ;
      RECT 128.78 22.25 129.04 22.57 ;
      RECT 128.84 19.87 128.98 22.57 ;
      RECT 128.78 19.87 129.04 20.19 ;
      RECT 126.02 29.39 126.28 29.71 ;
      RECT 126.02 29.48 126.68 29.62 ;
      RECT 126.54 24.04 126.68 29.62 ;
      RECT 126.08 24.04 126.68 24.18 ;
      RECT 126.08 22.59 126.22 24.18 ;
      RECT 126.02 22.59 126.28 22.91 ;
      RECT 126.02 16.13 126.28 16.45 ;
      RECT 126.08 11.37 126.22 16.45 ;
      RECT 126.02 11.37 126.28 11.69 ;
      RECT 126.02 30.41 126.28 30.73 ;
      RECT 125.62 30.5 126.28 30.64 ;
      RECT 125.62 16.9 125.76 30.64 ;
      RECT 126.02 16.81 126.28 17.13 ;
      RECT 125.62 16.9 126.28 17.04 ;
      RECT 126.02 21.23 126.28 21.55 ;
      RECT 126.08 17.49 126.22 21.55 ;
      RECT 126.02 17.49 126.28 17.81 ;
      RECT 126.02 26.67 126.28 26.99 ;
      RECT 126.08 24.63 126.22 26.99 ;
      RECT 126.02 24.63 126.28 24.95 ;
      RECT 123.26 13.41 123.52 13.73 ;
      RECT 123.32 12.05 123.46 13.73 ;
      RECT 123.26 12.05 123.52 12.37 ;
      RECT 123.26 16.13 123.52 16.45 ;
      RECT 123.32 14.77 123.46 16.45 ;
      RECT 123.26 14.77 123.52 15.09 ;
      RECT 123.26 18.51 123.52 18.83 ;
      RECT 123.32 17.15 123.46 18.83 ;
      RECT 123.26 17.15 123.52 17.47 ;
      RECT 123.26 32.11 123.52 32.43 ;
      RECT 123.32 28.03 123.46 32.43 ;
      RECT 123.26 30.07 123.52 30.39 ;
      RECT 123.26 28.03 123.52 28.35 ;
      RECT 122.86 28.12 123.52 28.26 ;
      RECT 122.86 21.32 123 28.26 ;
      RECT 122.86 21.32 123.46 21.46 ;
      RECT 123.32 19.19 123.46 21.46 ;
      RECT 123.26 19.19 123.52 19.51 ;
      RECT 123.26 27.35 123.52 27.67 ;
      RECT 123.32 22.25 123.46 27.67 ;
      RECT 123.26 22.25 123.52 22.57 ;
      RECT 120.5 18.85 120.76 19.17 ;
      RECT 120.56 17.24 120.7 19.17 ;
      RECT 120.1 17.24 120.7 17.38 ;
      RECT 120.1 13.84 120.24 17.38 ;
      RECT 120.1 13.84 120.7 13.98 ;
      RECT 120.56 13.07 120.7 13.98 ;
      RECT 120.5 13.07 120.76 13.39 ;
      RECT 120.5 30.07 120.76 30.39 ;
      RECT 120.56 27.01 120.7 30.39 ;
      RECT 120.5 27.69 120.76 28.01 ;
      RECT 120.5 27.01 120.76 27.33 ;
      RECT 118.14 16.13 118.4 16.45 ;
      RECT 118.2 14.43 118.34 16.45 ;
      RECT 118.14 14.43 118.4 14.75 ;
      RECT 117.74 13.75 118 14.07 ;
      RECT 117.8 12.05 117.94 14.07 ;
      RECT 117.74 12.05 118 12.37 ;
      RECT 117.74 18.85 118 19.17 ;
      RECT 117.8 16.81 117.94 19.17 ;
      RECT 117.74 16.81 118 17.13 ;
      RECT 117.74 24.63 118 24.95 ;
      RECT 117.8 19.53 117.94 24.95 ;
      RECT 117.74 22.25 118 22.57 ;
      RECT 117.74 19.53 118 19.85 ;
      RECT 117.74 38.23 118 38.55 ;
      RECT 117.8 25.65 117.94 38.55 ;
      RECT 117.74 28.03 118 28.35 ;
      RECT 117.74 25.65 118 25.97 ;
      RECT 114.98 18.51 115.24 18.83 ;
      RECT 115.04 14.865 115.18 18.83 ;
      RECT 114.97 14.865 115.25 15.235 ;
      RECT 114.98 29.39 115.24 29.71 ;
      RECT 115.04 19.19 115.18 29.71 ;
      RECT 114.98 21.23 115.24 21.55 ;
      RECT 114.98 19.19 115.24 19.51 ;
      RECT 112.19 27.04 112.51 27.3 ;
      RECT 111.82 27.1 112.51 27.24 ;
      RECT 111.82 24.72 111.96 27.24 ;
      RECT 111.82 24.72 112.42 24.86 ;
      RECT 112.28 23.36 112.42 24.86 ;
      RECT 112.22 23.95 112.48 24.27 ;
      RECT 112.28 23.36 112.88 23.5 ;
      RECT 112.74 15.88 112.88 23.5 ;
      RECT 112.22 16.81 112.48 17.13 ;
      RECT 112.28 15.79 112.42 17.13 ;
      RECT 112.22 15.79 112.48 16.11 ;
      RECT 112.22 15.88 112.88 16.02 ;
      RECT 112.22 32.11 112.48 32.43 ;
      RECT 112.22 32.2 112.88 32.34 ;
      RECT 112.74 26.76 112.88 32.34 ;
      RECT 112.22 30.75 112.48 31.07 ;
      RECT 112.22 30.84 112.88 30.98 ;
      RECT 112.28 26.76 112.88 26.9 ;
      RECT 112.28 25.65 112.42 26.9 ;
      RECT 112.22 25.65 112.48 25.97 ;
      RECT 112.21 14.865 112.49 15.235 ;
      RECT 112.28 13.75 112.42 15.235 ;
      RECT 112.22 13.75 112.48 14.07 ;
      RECT 112.22 22.59 112.48 22.91 ;
      RECT 112.28 21.66 112.42 22.91 ;
      RECT 112.05 21.66 112.42 21.8 ;
      RECT 112.05 18.6 112.19 21.8 ;
      RECT 112.05 18.6 112.42 18.74 ;
      RECT 112.28 17.49 112.42 18.74 ;
      RECT 112.22 17.49 112.48 17.81 ;
      RECT 112.22 30.07 112.48 30.39 ;
      RECT 112.28 27.69 112.42 30.39 ;
      RECT 112.22 27.69 112.48 28.01 ;
      RECT 109.46 27.69 109.72 28.01 ;
      RECT 109.52 16.56 109.66 28.01 ;
      RECT 109.46 24.63 109.72 24.95 ;
      RECT 109.46 17.49 109.72 17.81 ;
      RECT 109.52 16.56 110.12 16.7 ;
      RECT 109.98 14.52 110.12 16.7 ;
      RECT 109.43 14.46 109.75 14.72 ;
      RECT 109.43 14.52 110.12 14.66 ;
      RECT 109.46 15.79 109.72 16.11 ;
      RECT 109.52 14.865 109.66 16.11 ;
      RECT 109.45 14.865 109.73 15.235 ;
      RECT 109.45 30.115 109.73 30.485 ;
      RECT 109.52 29.39 109.66 30.485 ;
      RECT 109.46 29.39 109.72 29.71 ;
      RECT 103.94 17.49 104.2 17.81 ;
      RECT 104 15.79 104.14 17.81 ;
      RECT 103.94 15.79 104.2 16.11 ;
      RECT 101.18 21.23 101.44 21.55 ;
      RECT 101.24 16.81 101.38 21.55 ;
      RECT 101.18 16.81 101.44 17.13 ;
      RECT 101.18 29.39 101.44 29.71 ;
      RECT 101.24 22.59 101.38 29.71 ;
      RECT 101.18 22.59 101.44 22.91 ;
      RECT 98.42 28.03 98.68 28.35 ;
      RECT 98.48 11.37 98.62 28.35 ;
      RECT 98.42 23.95 98.68 24.27 ;
      RECT 98.42 13.07 98.68 13.39 ;
      RECT 98.42 11.37 98.68 11.69 ;
      RECT 95.66 23.95 95.92 24.27 ;
      RECT 95.72 22 95.86 24.27 ;
      RECT 95.72 22 96.32 22.14 ;
      RECT 96.18 13.16 96.32 22.14 ;
      RECT 95.66 13.07 95.92 13.39 ;
      RECT 95.66 13.16 96.32 13.3 ;
      RECT 95.65 30.115 95.93 30.485 ;
      RECT 95.66 30.07 95.92 30.485 ;
      RECT 95.66 18.85 95.92 19.17 ;
      RECT 95.72 13.75 95.86 19.17 ;
      RECT 95.66 16.81 95.92 17.13 ;
      RECT 95.66 13.75 95.92 14.07 ;
      RECT 95.66 29.39 95.92 29.71 ;
      RECT 95.72 24.72 95.86 29.71 ;
      RECT 95.26 24.72 95.86 24.86 ;
      RECT 95.26 21.32 95.4 24.86 ;
      RECT 95.26 21.32 95.86 21.46 ;
      RECT 95.72 20.21 95.86 21.46 ;
      RECT 95.66 20.21 95.92 20.53 ;
      RECT 92.9 16.47 93.16 16.79 ;
      RECT 92.96 13.07 93.1 16.79 ;
      RECT 92.89 14.865 93.17 15.235 ;
      RECT 92.9 13.07 93.16 13.39 ;
      RECT 92.89 30.725 93.17 31.095 ;
      RECT 92.96 27.69 93.1 31.095 ;
      RECT 92.9 29.73 93.16 30.05 ;
      RECT 92.9 27.69 93.16 28.01 ;
      RECT 92.9 18.85 93.16 19.17 ;
      RECT 92.96 17.49 93.1 19.17 ;
      RECT 92.9 17.49 93.16 17.81 ;
      RECT 92.9 22.25 93.16 22.57 ;
      RECT 92.96 19.53 93.1 22.57 ;
      RECT 92.9 19.53 93.16 19.85 ;
      RECT 92.9 27.01 93.16 27.33 ;
      RECT 92.96 22.93 93.1 27.33 ;
      RECT 92.9 22.93 93.16 23.25 ;
      RECT 90.14 21.23 90.4 21.55 ;
      RECT 90.2 11.37 90.34 21.55 ;
      RECT 90.14 18.85 90.4 19.17 ;
      RECT 90.14 14.43 90.4 14.75 ;
      RECT 90.14 11.37 90.4 11.69 ;
      RECT 90.14 24.63 90.4 24.95 ;
      RECT 90.2 22.25 90.34 24.95 ;
      RECT 90.14 22.25 90.4 22.57 ;
      RECT 90.14 29.73 90.4 30.05 ;
      RECT 90.2 28.37 90.34 30.05 ;
      RECT 90.14 28.37 90.4 28.69 ;
      RECT 87.38 18.51 87.64 18.83 ;
      RECT 87.38 18.6 88.04 18.74 ;
      RECT 87.9 11.8 88.04 18.74 ;
      RECT 87.38 11.71 87.64 12.03 ;
      RECT 87.38 11.8 88.04 11.94 ;
      RECT 87.38 16.81 87.64 17.13 ;
      RECT 87.44 14.77 87.58 17.13 ;
      RECT 87.38 15.79 87.64 16.11 ;
      RECT 87.38 14.77 87.64 15.09 ;
      RECT 87.38 31.09 87.64 31.41 ;
      RECT 87.44 19.53 87.58 31.41 ;
      RECT 87.38 19.53 87.64 19.85 ;
      RECT 84.62 16.13 84.88 16.45 ;
      RECT 84.68 14.865 84.82 16.45 ;
      RECT 84.61 14.865 84.89 15.235 ;
      RECT 84.62 23.95 84.88 24.27 ;
      RECT 84.68 22 84.82 24.27 ;
      RECT 84.22 22 84.82 22.14 ;
      RECT 84.22 18.6 84.36 22.14 ;
      RECT 84.62 18.51 84.88 18.83 ;
      RECT 84.22 18.6 84.88 18.74 ;
      RECT 84.62 21.23 84.88 21.55 ;
      RECT 84.68 20.21 84.82 21.55 ;
      RECT 84.62 20.21 84.88 20.53 ;
      RECT 84.62 29.39 84.88 29.71 ;
      RECT 84.68 27.35 84.82 29.71 ;
      RECT 84.62 27.35 84.88 27.67 ;
      RECT 84.62 32.11 84.88 32.43 ;
      RECT 84.68 30.41 84.82 32.43 ;
      RECT 84.62 30.41 84.88 30.73 ;
      RECT 81.92 20.64 82.52 20.78 ;
      RECT 82.38 14.98 82.52 20.78 ;
      RECT 81.92 19.53 82.06 20.78 ;
      RECT 81.86 19.53 82.12 19.85 ;
      RECT 82.305 13.75 82.445 15.12 ;
      RECT 82.245 13.75 82.505 14.07 ;
      RECT 81.85 25.845 82.13 26.215 ;
      RECT 81.92 22.93 82.06 26.215 ;
      RECT 81.86 22.93 82.12 23.25 ;
      RECT 81.86 16.13 82.12 16.45 ;
      RECT 81.92 11.37 82.06 16.45 ;
      RECT 81.86 11.37 82.12 11.69 ;
      RECT 81.86 18.85 82.12 19.17 ;
      RECT 81.92 17.49 82.06 19.17 ;
      RECT 81.86 17.49 82.12 17.81 ;
      RECT 81.86 32.11 82.12 32.43 ;
      RECT 81.92 30.75 82.06 32.43 ;
      RECT 81.86 30.75 82.12 31.07 ;
      RECT 79.1 20.21 79.36 20.53 ;
      RECT 78.7 20.3 79.36 20.44 ;
      RECT 78.7 15.88 78.84 20.44 ;
      RECT 79.1 16.81 79.36 17.13 ;
      RECT 79.16 14.865 79.3 17.13 ;
      RECT 78.7 15.88 79.3 16.02 ;
      RECT 79.09 14.865 79.37 15.235 ;
      RECT 79.09 30.115 79.37 30.485 ;
      RECT 79.1 30.07 79.36 30.485 ;
      RECT 79.1 18.85 79.36 19.17 ;
      RECT 79.16 17.49 79.3 19.17 ;
      RECT 79.1 17.49 79.36 17.81 ;
      RECT 79.1 29.39 79.36 29.71 ;
      RECT 79.16 24.29 79.3 29.71 ;
      RECT 79.1 24.29 79.36 24.61 ;
      RECT 76.34 29.39 76.6 29.71 ;
      RECT 76.4 17.915 76.54 29.71 ;
      RECT 76.34 22.93 76.6 23.25 ;
      RECT 76.33 17.915 76.61 18.285 ;
      RECT 76.34 32.45 76.6 32.77 ;
      RECT 76.4 30.07 76.54 32.77 ;
      RECT 76.34 31.09 76.6 31.41 ;
      RECT 76.34 30.07 76.6 30.39 ;
      RECT 73.58 32.11 73.84 32.43 ;
      RECT 73.64 30.75 73.78 32.43 ;
      RECT 73.58 30.75 73.84 31.07 ;
      RECT 73.58 30.84 74.24 30.98 ;
      RECT 74.1 16.56 74.24 30.98 ;
      RECT 73.58 27.01 73.84 27.33 ;
      RECT 73.58 27.1 74.24 27.24 ;
      RECT 73.58 16.47 73.84 16.79 ;
      RECT 73.58 16.56 74.24 16.7 ;
      RECT 73.58 11.37 73.84 11.69 ;
      RECT 73.64 10.595 73.78 11.69 ;
      RECT 73.57 10.595 73.85 10.965 ;
      RECT 73.57 25.845 73.85 26.215 ;
      RECT 73.64 19.19 73.78 26.215 ;
      RECT 73.58 24.97 73.84 25.29 ;
      RECT 73.58 19.19 73.84 19.51 ;
      RECT 73.57 30.115 73.85 30.485 ;
      RECT 73.18 30.16 73.85 30.3 ;
      RECT 73.18 27.78 73.32 30.3 ;
      RECT 73.58 30.07 73.84 30.485 ;
      RECT 73.58 27.69 73.84 28.01 ;
      RECT 73.18 27.78 73.84 27.92 ;
      RECT 73.58 15.79 73.84 16.11 ;
      RECT 73.64 13.07 73.78 16.11 ;
      RECT 73.58 13.07 73.84 13.39 ;
      RECT 73.58 18.51 73.84 18.83 ;
      RECT 73.64 17.49 73.78 18.83 ;
      RECT 73.58 17.49 73.84 17.81 ;
      RECT 73.58 29.39 73.84 29.71 ;
      RECT 73.64 28.37 73.78 29.71 ;
      RECT 73.58 28.37 73.84 28.69 ;
      RECT 70.82 31.09 71.08 31.41 ;
      RECT 70.88 18.6 71.02 31.41 ;
      RECT 70.88 18.6 71.48 18.74 ;
      RECT 71.34 17.92 71.48 18.74 ;
      RECT 70.88 17.92 71.48 18.06 ;
      RECT 70.88 17.52 71.02 18.06 ;
      RECT 70.79 17.52 71.11 17.78 ;
      RECT 70.82 16.13 71.08 16.45 ;
      RECT 70.88 13.75 71.02 16.45 ;
      RECT 70.82 13.75 71.08 14.07 ;
      RECT 68.06 23.95 68.32 24.27 ;
      RECT 68.06 24.04 68.72 24.18 ;
      RECT 68.58 16.56 68.72 24.18 ;
      RECT 68.06 16.47 68.32 16.79 ;
      RECT 68.06 16.56 68.72 16.7 ;
      RECT 68.12 14.77 68.26 16.79 ;
      RECT 68.06 14.77 68.32 15.09 ;
      RECT 68.06 27.69 68.32 28.01 ;
      RECT 68.12 24.72 68.26 28.01 ;
      RECT 67.66 24.72 68.26 24.86 ;
      RECT 67.66 23.02 67.8 24.86 ;
      RECT 67.66 23.02 68.03 23.16 ;
      RECT 67.89 18.6 68.03 23.16 ;
      RECT 67.89 18.6 68.26 18.74 ;
      RECT 68.12 17.49 68.26 18.74 ;
      RECT 68.06 17.49 68.32 17.81 ;
      RECT 65.29 25.845 65.57 26.215 ;
      RECT 65.36 22.25 65.5 26.215 ;
      RECT 65.3 22.25 65.56 22.57 ;
      RECT 65.3 32.45 65.56 32.77 ;
      RECT 65.36 27.065 65.5 32.77 ;
      RECT 65.3 27.065 65.56 27.67 ;
      RECT 65.29 27.065 65.57 27.435 ;
      RECT 65.3 19.53 65.56 19.85 ;
      RECT 65.36 12.05 65.5 19.85 ;
      RECT 65.3 15.79 65.56 16.11 ;
      RECT 65.3 12.05 65.56 12.37 ;
      RECT 62.54 18.51 62.8 18.83 ;
      RECT 62.54 18.6 63.2 18.74 ;
      RECT 63.06 13.84 63.2 18.74 ;
      RECT 62.54 13.645 62.8 14.07 ;
      RECT 62.53 13.645 62.81 14.015 ;
      RECT 62.53 13.84 63.2 13.98 ;
      RECT 62.54 21.23 62.8 21.55 ;
      RECT 62.6 19.28 62.74 21.55 ;
      RECT 62.14 19.28 62.74 19.42 ;
      RECT 62.14 13.16 62.28 19.42 ;
      RECT 62.54 13.07 62.8 13.39 ;
      RECT 62.14 13.16 62.8 13.3 ;
      RECT 62.6 11.37 62.74 13.39 ;
      RECT 62.54 11.37 62.8 11.69 ;
      RECT 62.54 16.81 62.8 17.13 ;
      RECT 62.6 14.77 62.74 17.13 ;
      RECT 62.54 14.77 62.8 15.09 ;
      RECT 62.54 26.67 62.8 26.99 ;
      RECT 62.6 25.31 62.74 26.99 ;
      RECT 62.54 25.31 62.8 25.63 ;
      RECT 62.54 29.73 62.8 30.05 ;
      RECT 62.6 28.37 62.74 30.05 ;
      RECT 62.54 28.37 62.8 28.69 ;
      RECT 59.77 14.865 60.05 15.235 ;
      RECT 59.84 14.09 59.98 15.235 ;
      RECT 59.78 14.09 60.04 14.41 ;
      RECT 59.78 30.07 60.04 30.39 ;
      RECT 59.84 16.81 59.98 30.39 ;
      RECT 59.78 27.69 60.04 28.01 ;
      RECT 59.78 22.795 60.04 23.25 ;
      RECT 59.77 22.795 60.05 23.165 ;
      RECT 59.78 19.19 60.04 19.51 ;
      RECT 59.78 16.81 60.04 17.13 ;
      RECT 57.02 21.23 57.28 21.55 ;
      RECT 56.62 21.32 57.28 21.46 ;
      RECT 56.62 13.84 56.76 21.46 ;
      RECT 57.02 18.51 57.28 18.83 ;
      RECT 56.62 18.6 57.28 18.74 ;
      RECT 57.02 17.15 57.28 17.47 ;
      RECT 56.62 17.24 57.28 17.38 ;
      RECT 57.02 13.75 57.28 14.07 ;
      RECT 56.62 13.84 57.28 13.98 ;
      RECT 57.02 32.11 57.28 32.43 ;
      RECT 57.08 28.03 57.22 32.43 ;
      RECT 57.02 28.03 57.28 28.35 ;
      RECT 54.26 30.07 54.52 30.39 ;
      RECT 54.32 27.065 54.46 30.39 ;
      RECT 54.26 27.065 54.52 27.67 ;
      RECT 54.25 27.065 54.53 27.435 ;
      RECT 54.26 18.85 54.52 19.17 ;
      RECT 54.32 14.77 54.46 19.17 ;
      RECT 54.26 14.77 54.52 15.09 ;
      RECT 54.26 22.59 54.52 22.91 ;
      RECT 54.32 20.21 54.46 22.91 ;
      RECT 54.26 20.21 54.52 20.53 ;
      RECT 54.26 34.83 54.52 35.15 ;
      RECT 54.32 30.75 54.46 35.15 ;
      RECT 54.26 30.75 54.52 31.07 ;
      RECT 51.5 27.35 51.76 27.67 ;
      RECT 51.56 25.4 51.7 27.67 ;
      RECT 51.56 25.4 52.16 25.54 ;
      RECT 52.02 22 52.16 25.54 ;
      RECT 51.56 22 52.16 22.14 ;
      RECT 51.56 21.23 51.7 22.14 ;
      RECT 51.5 21.23 51.76 21.55 ;
      RECT 51.5 35.17 51.76 35.49 ;
      RECT 51.56 34.24 51.7 35.49 ;
      RECT 51.56 34.24 52.16 34.38 ;
      RECT 52.02 30.16 52.16 34.38 ;
      RECT 51.56 30.16 52.16 30.3 ;
      RECT 51.56 28.37 51.7 30.3 ;
      RECT 51.5 28.37 51.76 28.69 ;
      RECT 51.49 14.255 51.77 14.625 ;
      RECT 51.5 14.09 51.76 14.625 ;
      RECT 51.5 13.07 51.76 13.39 ;
      RECT 51.56 12.05 51.7 13.39 ;
      RECT 51.5 12.05 51.76 12.37 ;
      RECT 51.5 16.81 51.76 17.13 ;
      RECT 51.56 14.77 51.7 17.13 ;
      RECT 51.5 14.77 51.76 15.09 ;
      RECT 51.5 18.85 51.76 19.17 ;
      RECT 51.56 17.49 51.7 19.17 ;
      RECT 51.5 17.49 51.76 17.81 ;
      RECT 51.5 24.29 51.76 24.61 ;
      RECT 51.56 22.93 51.7 24.61 ;
      RECT 51.5 22.93 51.76 23.25 ;
      RECT 51.5 33.13 51.76 33.45 ;
      RECT 51.56 31.09 51.7 33.45 ;
      RECT 51.5 31.09 51.76 31.41 ;
      RECT 48.74 15.79 49 16.11 ;
      RECT 48.8 13.84 48.94 16.11 ;
      RECT 48.8 13.84 49.4 13.98 ;
      RECT 49.26 11.8 49.4 13.98 ;
      RECT 48.34 11.8 49.4 11.94 ;
      RECT 48.34 9.33 48.48 11.94 ;
      RECT 48.28 9.33 48.54 9.65 ;
      RECT 48.395 18.51 48.655 18.83 ;
      RECT 48.455 17.92 48.595 18.83 ;
      RECT 48.34 13.16 48.48 18.06 ;
      RECT 48.34 14.43 48.655 14.75 ;
      RECT 48.71 13.44 49.03 13.7 ;
      RECT 48.8 13.16 48.94 13.7 ;
      RECT 48.34 13.16 48.94 13.3 ;
      RECT 48.74 35.51 49 35.83 ;
      RECT 48.8 16.81 48.94 35.83 ;
      RECT 48.74 32.79 49 33.11 ;
      RECT 48.74 24.63 49 24.95 ;
      RECT 48.73 22.795 49.01 23.165 ;
      RECT 48.74 19.19 49 19.51 ;
      RECT 48.74 16.81 49 17.13 ;
      RECT 45.98 15.79 46.24 16.11 ;
      RECT 45.98 15.88 46.64 16.02 ;
      RECT 46.5 8.765 46.64 16.02 ;
      RECT 45.98 13.07 46.24 13.39 ;
      RECT 45.98 13.16 46.64 13.3 ;
      RECT 46.43 8.765 46.71 9.135 ;
      RECT 45.98 30.07 46.24 30.39 ;
      RECT 46.04 27.69 46.18 30.39 ;
      RECT 45.98 29.39 46.24 29.71 ;
      RECT 46.04 28.8 46.64 28.94 ;
      RECT 46.5 21.32 46.64 28.94 ;
      RECT 45.98 27.69 46.24 28.01 ;
      RECT 45.98 22.25 46.24 22.57 ;
      RECT 46.04 16.47 46.18 22.57 ;
      RECT 46.04 21.32 46.64 21.46 ;
      RECT 45.98 16.47 46.24 16.79 ;
      RECT 45.98 26.67 46.24 26.99 ;
      RECT 46.04 24.32 46.18 26.99 ;
      RECT 45.95 24.32 46.27 24.58 ;
      RECT 45.98 14.43 46.24 14.75 ;
      RECT 45.58 14.52 46.24 14.66 ;
      RECT 45.58 12.48 45.72 14.66 ;
      RECT 45.58 12.48 46.18 12.62 ;
      RECT 46.04 11.37 46.18 12.62 ;
      RECT 45.98 11.37 46.24 11.69 ;
      RECT 45.98 30.75 46.24 31.07 ;
      RECT 45.58 30.84 46.24 30.98 ;
      RECT 45.58 24.04 45.72 30.98 ;
      RECT 45.58 24.04 46.18 24.18 ;
      RECT 46.04 22.93 46.18 24.18 ;
      RECT 45.98 22.93 46.24 23.25 ;
      RECT 43.22 30.41 43.48 30.73 ;
      RECT 43.28 16.56 43.42 30.73 ;
      RECT 43.22 27.35 43.48 27.67 ;
      RECT 43.22 21.91 43.48 22.23 ;
      RECT 43.22 17.15 43.48 17.47 ;
      RECT 43.28 16.56 43.88 16.7 ;
      RECT 43.74 13.84 43.88 16.7 ;
      RECT 43.28 13.84 43.88 13.98 ;
      RECT 43.28 13.44 43.42 13.98 ;
      RECT 43.19 13.44 43.51 13.7 ;
      RECT 43.19 14.12 43.51 14.38 ;
      RECT 42.82 14.18 43.51 14.32 ;
      RECT 42.82 9.33 42.96 14.32 ;
      RECT 42.76 9.33 43.02 9.65 ;
      RECT 43.19 16.16 43.51 16.42 ;
      RECT 43.28 14.77 43.42 16.42 ;
      RECT 43.21 14.865 43.49 15.235 ;
      RECT 43.22 14.77 43.48 15.235 ;
      RECT 40.46 38.23 40.72 38.55 ;
      RECT 40.52 30.84 40.66 38.55 ;
      RECT 40.52 30.84 41.12 30.98 ;
      RECT 40.98 22.68 41.12 30.98 ;
      RECT 40.46 22.59 40.72 22.91 ;
      RECT 40.46 22.68 41.12 22.82 ;
      RECT 40.46 29.73 40.72 30.05 ;
      RECT 40.52 28.8 40.66 30.05 ;
      RECT 40.29 28.8 40.66 28.94 ;
      RECT 40.29 23.7 40.43 28.94 ;
      RECT 40.06 23.7 40.43 23.84 ;
      RECT 40.06 22 40.2 23.84 ;
      RECT 40.06 22 40.66 22.14 ;
      RECT 40.52 16.81 40.66 22.14 ;
      RECT 40.46 16.81 40.72 17.13 ;
      RECT 34.94 17.49 35.2 17.81 ;
      RECT 35 14.77 35.14 17.81 ;
      RECT 34.94 14.77 35.2 15.09 ;
      RECT 32.18 21.23 32.44 21.55 ;
      RECT 32.24 17.15 32.38 21.55 ;
      RECT 32.18 17.15 32.44 17.47 ;
      RECT 29.42 22.59 29.68 22.91 ;
      RECT 29.48 17.15 29.62 22.91 ;
      RECT 29.42 17.15 29.68 17.47 ;
    LAYER via2 ;
      RECT 170.21 18.61 170.41 18.81 ;
      RECT 164.69 18.61 164.89 18.81 ;
      RECT 164.69 25.93 164.89 26.13 ;
      RECT 161.93 18.61 162.13 18.81 ;
      RECT 153.65 18.61 153.85 18.81 ;
      RECT 150.43 9.46 150.63 9.66 ;
      RECT 142.61 14.95 142.81 15.15 ;
      RECT 142.61 18.61 142.81 18.81 ;
      RECT 140.31 9.46 140.51 9.66 ;
      RECT 131.57 14.95 131.77 15.15 ;
      RECT 131.57 25.93 131.77 26.13 ;
      RECT 128.81 18 129.01 18.2 ;
      RECT 115.01 14.95 115.21 15.15 ;
      RECT 112.25 14.95 112.45 15.15 ;
      RECT 109.49 14.95 109.69 15.15 ;
      RECT 109.49 30.2 109.69 30.4 ;
      RECT 95.69 30.2 95.89 30.4 ;
      RECT 92.93 14.95 93.13 15.15 ;
      RECT 92.93 30.81 93.13 31.01 ;
      RECT 84.65 14.95 84.85 15.15 ;
      RECT 81.89 25.93 82.09 26.13 ;
      RECT 79.13 14.95 79.33 15.15 ;
      RECT 79.13 30.2 79.33 30.4 ;
      RECT 76.37 18 76.57 18.2 ;
      RECT 73.61 10.68 73.81 10.88 ;
      RECT 73.61 25.93 73.81 26.13 ;
      RECT 73.61 30.2 73.81 30.4 ;
      RECT 65.33 25.93 65.53 26.13 ;
      RECT 65.33 27.15 65.53 27.35 ;
      RECT 62.57 13.73 62.77 13.93 ;
      RECT 59.81 14.95 60.01 15.15 ;
      RECT 59.81 22.88 60.01 23.08 ;
      RECT 54.29 27.15 54.49 27.35 ;
      RECT 51.53 14.34 51.73 14.54 ;
      RECT 48.77 22.88 48.97 23.08 ;
      RECT 46.47 8.85 46.67 9.05 ;
      RECT 43.25 14.95 43.45 15.15 ;
    LAYER met3 ;
      RECT 170.145 18.545 170.475 18.875 ;
      RECT 164.625 18.545 164.955 18.875 ;
      RECT 161.865 18.545 162.195 18.875 ;
      RECT 153.585 18.545 153.915 18.875 ;
      RECT 153.585 18.56 170.475 18.86 ;
      RECT 132.9 26.49 163.56 26.79 ;
      RECT 163.26 25.88 163.56 26.79 ;
      RECT 132.9 25.88 133.2 26.79 ;
      RECT 164.625 25.865 164.955 26.195 ;
      RECT 131.505 25.865 131.835 26.195 ;
      RECT 163.26 25.88 164.955 26.18 ;
      RECT 131.505 25.88 133.2 26.18 ;
      RECT 150.365 9.395 150.695 9.725 ;
      RECT 140.245 9.395 140.575 9.725 ;
      RECT 140.245 9.41 150.695 9.71 ;
      RECT 142.545 14.885 142.875 15.215 ;
      RECT 131.505 14.885 131.835 15.215 ;
      RECT 141.18 14.9 142.875 15.2 ;
      RECT 131.505 14.9 133.2 15.2 ;
      RECT 132.9 14.29 133.2 15.2 ;
      RECT 141.18 14.29 141.48 15.2 ;
      RECT 132.9 14.29 141.48 14.59 ;
      RECT 142.545 18.545 142.875 18.875 ;
      RECT 138.42 18.56 142.875 18.86 ;
      RECT 138.42 18.255 138.72 18.86 ;
      RECT 130.14 18.255 138.72 18.555 ;
      RECT 128.745 17.935 129.075 18.265 ;
      RECT 130.14 17.95 130.44 18.555 ;
      RECT 128.745 17.95 130.44 18.25 ;
      RECT 114.945 14.885 115.275 15.215 ;
      RECT 112.185 14.885 112.515 15.215 ;
      RECT 112.185 14.9 115.275 15.2 ;
      RECT 109.425 14.885 109.755 15.215 ;
      RECT 92.865 14.885 93.195 15.215 ;
      RECT 108.06 14.9 109.755 15.2 ;
      RECT 92.865 14.9 94.56 15.2 ;
      RECT 94.26 14.29 94.56 15.2 ;
      RECT 108.06 14.29 108.36 15.2 ;
      RECT 94.26 14.29 108.36 14.59 ;
      RECT 97.02 30.455 108.36 30.755 ;
      RECT 108.06 30.15 108.36 30.755 ;
      RECT 109.425 30.135 109.755 30.465 ;
      RECT 95.625 30.135 95.955 30.465 ;
      RECT 97.02 30.15 97.32 30.755 ;
      RECT 108.06 30.15 109.755 30.45 ;
      RECT 95.625 30.15 97.32 30.45 ;
      RECT 92.865 30.745 93.195 31.075 ;
      RECT 86.9 30.76 93.195 31.06 ;
      RECT 86.9 30.455 87.2 31.06 ;
      RECT 80.46 30.455 87.2 30.755 ;
      RECT 79.065 30.135 79.395 30.465 ;
      RECT 73.545 30.135 73.875 30.465 ;
      RECT 80.46 30.15 80.76 30.755 ;
      RECT 73.545 30.15 80.76 30.45 ;
      RECT 84.585 14.885 84.915 15.215 ;
      RECT 79.065 14.885 79.395 15.215 ;
      RECT 59.745 14.885 60.075 15.215 ;
      RECT 77.7 14.9 84.915 15.2 ;
      RECT 59.745 14.9 64.2 15.2 ;
      RECT 63.9 14.29 64.2 15.2 ;
      RECT 77.7 14.29 78 15.2 ;
      RECT 63.9 14.29 78 14.59 ;
      RECT 81.825 25.865 82.155 26.195 ;
      RECT 73.545 25.865 73.875 26.195 ;
      RECT 65.265 25.865 65.595 26.195 ;
      RECT 65.265 25.88 82.155 26.18 ;
      RECT 73.545 10.615 73.875 10.945 ;
      RECT 76.28 10.62 76.66 10.94 ;
      RECT 73.545 10.63 76.66 10.93 ;
      RECT 76.305 17.935 76.635 18.265 ;
      RECT 76.28 17.94 76.66 18.26 ;
      RECT 75.86 17.95 76.66 18.25 ;
      RECT 65.265 27.085 65.595 27.415 ;
      RECT 54.225 27.085 54.555 27.415 ;
      RECT 63.9 27.1 65.595 27.4 ;
      RECT 54.225 27.1 55.92 27.4 ;
      RECT 55.62 26.49 55.92 27.4 ;
      RECT 63.9 26.49 64.2 27.4 ;
      RECT 55.62 26.49 64.2 26.79 ;
      RECT 62.505 13.665 62.835 13.995 ;
      RECT 60.41 13.67 60.79 13.99 ;
      RECT 60.41 13.68 62.835 13.98 ;
      RECT 46.405 8.785 46.735 9.115 ;
      RECT 60.41 8.79 60.79 9.11 ;
      RECT 46.405 8.8 60.79 9.1 ;
      RECT 59.745 22.815 60.075 23.145 ;
      RECT 48.705 22.815 49.035 23.145 ;
      RECT 48.705 22.83 60.075 23.13 ;
      RECT 43.185 14.885 43.515 15.215 ;
      RECT 43.185 14.9 44.88 15.2 ;
      RECT 44.58 14.29 44.88 15.2 ;
      RECT 51.465 14.275 51.795 14.605 ;
      RECT 44.58 14.29 51.795 14.59 ;
    LAYER via3 ;
      RECT 76.37 10.68 76.57 10.88 ;
      RECT 76.37 18 76.57 18.2 ;
      RECT 60.5 8.85 60.7 9.05 ;
      RECT 60.5 13.73 60.7 13.93 ;
    LAYER met4 ;
      RECT 76.305 17.935 76.635 18.265 ;
      RECT 76.32 10.615 76.62 18.265 ;
      RECT 76.305 10.615 76.635 10.945 ;
      RECT 60.435 13.665 60.765 13.995 ;
      RECT 60.45 8.785 60.75 13.995 ;
      RECT 60.435 8.785 60.765 9.115 ;
    LAYER li1 ;
      RECT 183.875 22.775 184.205 23.295 ;
      RECT 184.085 22.025 184.255 22.86 ;
      RECT 184.03 22.735 184.255 22.86 ;
      RECT 184.04 22.025 184.255 22.155 ;
      RECT 183.865 21.18 184.195 22.105 ;
      RECT 181.135 25.045 181.465 26.065 ;
      RECT 180.295 25.045 180.625 26.065 ;
      RECT 180.295 25.045 181.795 25.215 ;
      RECT 181.62 24.335 181.795 25.215 ;
      RECT 181.62 24.675 184.245 24.845 ;
      RECT 180.375 24.335 181.795 24.505 ;
      RECT 181.215 23.86 181.385 24.505 ;
      RECT 180.375 23.855 180.545 24.505 ;
      RECT 183.035 22.775 183.365 23.3 ;
      RECT 183.165 22.275 183.365 23.3 ;
      RECT 183.165 22.275 183.915 22.605 ;
      RECT 183.165 21.135 183.355 23.3 ;
      RECT 182.46 21.695 183.355 22.07 ;
      RECT 183.015 21.135 183.355 22.07 ;
      RECT 181.505 23.065 182.29 23.235 ;
      RECT 182.12 21.265 182.29 23.235 ;
      RECT 182.12 22.275 182.995 22.605 ;
      RECT 181.405 21.265 182.29 21.435 ;
      RECT 181.485 22.565 181.95 22.895 ;
      RECT 181.63 21.605 181.95 22.895 ;
      RECT 180.93 23.065 181.335 23.235 ;
      RECT 180.93 21.135 181.1 23.235 ;
      RECT 180.27 22.535 181.1 22.835 ;
      RECT 180.27 22.505 180.47 22.835 ;
      RECT 180.93 21.135 181.18 21.465 ;
      RECT 177.155 17.255 177.325 17.905 ;
      RECT 177.995 17.255 178.165 17.9 ;
      RECT 177.155 17.255 178.575 17.425 ;
      RECT 178.4 16.545 178.575 17.425 ;
      RECT 178.4 16.915 181.025 17.085 ;
      RECT 177.075 16.545 178.575 16.715 ;
      RECT 177.915 15.695 178.245 16.715 ;
      RECT 177.075 15.695 177.405 16.715 ;
      RECT 179.385 23.065 180.06 23.235 ;
      RECT 179.89 22.115 180.06 23.235 ;
      RECT 180.59 22.025 180.76 22.355 ;
      RECT 179.89 22.115 180.76 22.285 ;
      RECT 180.25 22.025 180.76 22.285 ;
      RECT 180.25 21.24 180.42 22.285 ;
      RECT 179.315 21.24 180.42 21.41 ;
      RECT 179.195 22.645 179.72 22.865 ;
      RECT 179.55 21.58 179.72 22.865 ;
      RECT 179.55 21.58 180.08 21.945 ;
      RECT 178.855 23.065 179.19 23.235 ;
      RECT 178.855 22.795 179.025 23.235 ;
      RECT 178.8 21.56 178.97 22.925 ;
      RECT 178.855 21.135 179.105 21.69 ;
      RECT 177.155 22.795 177.325 23.255 ;
      RECT 177.155 22.795 177.82 22.965 ;
      RECT 177.59 21.635 177.82 22.965 ;
      RECT 177.155 21.635 177.82 21.805 ;
      RECT 177.155 21.135 177.325 21.805 ;
      RECT 176.055 17.335 176.385 17.855 ;
      RECT 176.265 16.585 176.435 17.42 ;
      RECT 176.21 17.295 176.435 17.42 ;
      RECT 176.22 16.585 176.435 16.715 ;
      RECT 176.045 15.74 176.375 16.665 ;
      RECT 175.215 17.335 175.545 17.86 ;
      RECT 175.345 16.835 175.545 17.86 ;
      RECT 175.345 16.835 176.095 17.165 ;
      RECT 175.345 15.695 175.535 17.86 ;
      RECT 174.64 16.255 175.535 16.63 ;
      RECT 175.195 15.695 175.535 16.63 ;
      RECT 173.685 17.625 174.47 17.795 ;
      RECT 174.3 15.825 174.47 17.795 ;
      RECT 174.3 16.835 175.175 17.165 ;
      RECT 173.585 15.825 174.47 15.995 ;
      RECT 173.9 20.015 174.085 20.595 ;
      RECT 173.9 20.015 174.565 20.19 ;
      RECT 174.225 18.815 174.565 20.19 ;
      RECT 173.88 18.815 174.565 18.985 ;
      RECT 173.88 18.415 174.085 18.985 ;
      RECT 173.665 17.125 174.13 17.455 ;
      RECT 173.81 16.165 174.13 17.455 ;
      RECT 172.925 19.655 173.195 20.595 ;
      RECT 172.925 19.655 174.055 19.825 ;
      RECT 173.805 19.155 174.055 19.825 ;
      RECT 172.925 18.415 173.095 20.595 ;
      RECT 172.925 18.415 173.185 18.745 ;
      RECT 173.11 17.625 173.515 17.795 ;
      RECT 173.11 15.695 173.28 17.795 ;
      RECT 172.45 17.095 173.28 17.395 ;
      RECT 172.45 17.065 172.65 17.395 ;
      RECT 173.11 15.695 173.36 16.025 ;
      RECT 172.5 22.775 172.705 23.345 ;
      RECT 172.5 22.775 173.185 22.945 ;
      RECT 172.845 21.57 173.185 22.945 ;
      RECT 172.52 21.57 173.185 21.745 ;
      RECT 172.52 21.165 172.705 21.745 ;
      RECT 171.565 17.625 172.24 17.795 ;
      RECT 172.07 16.675 172.24 17.795 ;
      RECT 172.77 16.585 172.94 16.915 ;
      RECT 172.07 16.675 172.94 16.845 ;
      RECT 172.43 16.585 172.94 16.845 ;
      RECT 172.43 15.8 172.6 16.845 ;
      RECT 171.495 15.8 172.6 15.97 ;
      RECT 172.365 19.655 172.695 20.58 ;
      RECT 172.585 18.9 172.755 19.735 ;
      RECT 172.54 19.605 172.755 19.735 ;
      RECT 172.53 18.9 172.755 19.025 ;
      RECT 172.375 18.465 172.705 18.985 ;
      RECT 171.545 23.015 171.805 23.345 ;
      RECT 171.545 21.165 171.715 23.345 ;
      RECT 172.425 21.935 172.675 22.605 ;
      RECT 171.545 21.935 172.675 22.105 ;
      RECT 171.545 21.165 171.815 22.105 ;
      RECT 171.515 19.69 171.855 20.625 ;
      RECT 171.665 18.46 171.855 20.625 ;
      RECT 170.96 19.69 171.855 20.065 ;
      RECT 171.665 19.155 172.415 19.485 ;
      RECT 171.665 18.46 171.865 19.485 ;
      RECT 171.535 18.46 171.865 18.985 ;
      RECT 171.375 17.205 171.9 17.425 ;
      RECT 171.73 16.14 171.9 17.425 ;
      RECT 171.73 16.14 172.26 16.505 ;
      RECT 171.555 25.105 171.815 26.055 ;
      RECT 170.655 25.105 170.885 26.055 ;
      RECT 170.655 25.105 171.815 25.345 ;
      RECT 169.905 20.325 170.79 20.495 ;
      RECT 170.62 18.525 170.79 20.495 ;
      RECT 170.62 19.155 171.495 19.485 ;
      RECT 170.005 18.525 170.79 18.695 ;
      RECT 171.115 22.84 171.375 23.345 ;
      RECT 171.205 21.135 171.375 23.345 ;
      RECT 171.105 21.135 171.375 22.04 ;
      RECT 171.035 17.625 171.37 17.795 ;
      RECT 171.035 17.355 171.205 17.795 ;
      RECT 170.98 16.12 171.15 17.485 ;
      RECT 171.035 15.695 171.285 16.25 ;
      RECT 170.82 24.615 171.345 24.925 ;
      RECT 171.115 23.975 171.345 24.925 ;
      RECT 171.115 14.175 171.285 15.185 ;
      RECT 168.225 14.175 171.285 14.345 ;
      RECT 168.225 13.455 168.395 14.345 ;
      RECT 170.22 13.455 171.285 13.625 ;
      RECT 171.115 12.975 171.285 13.625 ;
      RECT 168.225 13.455 169.025 13.625 ;
      RECT 168.855 12.975 169.025 13.625 ;
      RECT 170.22 12.975 170.39 13.625 ;
      RECT 168.855 12.975 170.39 13.225 ;
      RECT 170.255 22.795 170.425 23.345 ;
      RECT 170.255 22.795 170.92 22.965 ;
      RECT 170.75 21.895 170.92 22.965 ;
      RECT 170.75 22.21 171.035 22.54 ;
      RECT 170.255 21.895 170.92 22.065 ;
      RECT 170.255 21.135 170.425 22.065 ;
      RECT 169.775 15.015 170.945 15.185 ;
      RECT 170.615 14.515 170.945 15.185 ;
      RECT 169.775 14.975 170.105 15.185 ;
      RECT 170.205 25.105 170.475 26.055 ;
      RECT 169.705 25.105 170.475 25.325 ;
      RECT 169.705 24.235 169.995 25.325 ;
      RECT 169.705 24.235 170.935 24.435 ;
      RECT 170.625 23.865 170.935 24.435 ;
      RECT 170.13 18.865 170.45 20.155 ;
      RECT 169.985 18.865 170.45 19.195 ;
      RECT 168.81 14.515 169.06 15.185 ;
      RECT 170.215 14.515 170.445 14.845 ;
      RECT 168.81 14.515 170.445 14.755 ;
      RECT 169.76 13.795 170.235 13.995 ;
      RECT 169.76 13.395 170.04 13.995 ;
      RECT 169.335 17.355 169.505 17.815 ;
      RECT 169.335 17.355 170 17.525 ;
      RECT 169.77 16.195 170 17.525 ;
      RECT 169.335 16.195 170 16.365 ;
      RECT 169.335 15.695 169.505 16.365 ;
      RECT 169.43 20.295 169.68 20.625 ;
      RECT 169.43 18.525 169.6 20.625 ;
      RECT 168.77 18.925 168.97 19.255 ;
      RECT 168.77 18.925 169.6 19.225 ;
      RECT 169.43 18.525 169.835 18.695 ;
      RECT 169.155 22.775 169.485 23.295 ;
      RECT 169.365 22.025 169.535 22.86 ;
      RECT 169.31 22.735 169.535 22.86 ;
      RECT 169.32 22.025 169.535 22.155 ;
      RECT 169.145 21.18 169.475 22.105 ;
      RECT 169.16 13.795 169.49 13.995 ;
      RECT 169.205 13.395 169.49 13.995 ;
      RECT 167.815 20.35 168.92 20.52 ;
      RECT 168.75 19.475 168.92 20.52 ;
      RECT 168.75 19.475 169.26 19.735 ;
      RECT 169.09 19.405 169.26 19.735 ;
      RECT 168.39 19.475 169.26 19.645 ;
      RECT 168.39 18.525 168.56 19.645 ;
      RECT 167.885 18.525 168.56 18.695 ;
      RECT 168.315 22.775 168.645 23.3 ;
      RECT 168.445 22.275 168.645 23.3 ;
      RECT 168.445 22.275 169.195 22.605 ;
      RECT 168.445 21.135 168.635 23.3 ;
      RECT 167.74 21.695 168.635 22.07 ;
      RECT 168.295 21.135 168.635 22.07 ;
      RECT 168.615 13.825 168.99 13.995 ;
      RECT 168.625 13.795 168.99 13.995 ;
      RECT 168.05 19.815 168.58 20.18 ;
      RECT 168.05 18.895 168.22 20.18 ;
      RECT 167.695 18.895 168.22 19.115 ;
      RECT 166.785 23.065 167.57 23.235 ;
      RECT 167.4 21.265 167.57 23.235 ;
      RECT 167.4 22.275 168.275 22.605 ;
      RECT 166.685 21.265 167.57 21.435 ;
      RECT 167.885 14.515 168.14 15.185 ;
      RECT 167.885 12.975 168.055 15.185 ;
      RECT 167.885 12.975 168.07 13.385 ;
      RECT 167.885 12.975 168.14 13.305 ;
      RECT 167.355 20.07 167.605 20.625 ;
      RECT 167.3 18.835 167.47 20.2 ;
      RECT 167.355 18.525 167.525 18.965 ;
      RECT 167.355 18.525 167.69 18.695 ;
      RECT 166.765 22.565 167.23 22.895 ;
      RECT 166.91 21.605 167.23 22.895 ;
      RECT 163.355 11.815 163.525 12.465 ;
      RECT 164.195 11.815 164.365 12.46 ;
      RECT 163.355 11.815 164.775 11.985 ;
      RECT 164.6 11.105 164.775 11.985 ;
      RECT 164.6 11.475 167.225 11.645 ;
      RECT 163.275 11.105 164.775 11.275 ;
      RECT 164.115 10.255 164.445 11.275 ;
      RECT 163.275 10.255 163.605 11.275 ;
      RECT 166.21 23.065 166.615 23.235 ;
      RECT 166.21 21.135 166.38 23.235 ;
      RECT 165.55 22.535 166.38 22.835 ;
      RECT 165.55 22.505 165.75 22.835 ;
      RECT 166.21 21.135 166.46 21.465 ;
      RECT 165.655 19.955 165.825 20.625 ;
      RECT 165.655 19.955 166.32 20.125 ;
      RECT 166.09 18.795 166.32 20.125 ;
      RECT 165.655 18.795 166.32 18.965 ;
      RECT 165.655 18.505 165.825 18.965 ;
      RECT 162.435 17.255 162.605 17.905 ;
      RECT 163.275 17.255 163.445 17.9 ;
      RECT 162.435 17.255 163.855 17.425 ;
      RECT 163.68 16.545 163.855 17.425 ;
      RECT 163.68 16.915 166.305 17.085 ;
      RECT 162.355 16.545 163.855 16.715 ;
      RECT 163.195 15.695 163.525 16.715 ;
      RECT 162.355 15.695 162.685 16.715 ;
      RECT 164.665 23.065 165.34 23.235 ;
      RECT 165.17 22.115 165.34 23.235 ;
      RECT 165.87 22.025 166.04 22.355 ;
      RECT 165.17 22.115 166.04 22.285 ;
      RECT 165.53 22.025 166.04 22.285 ;
      RECT 165.53 21.24 165.7 22.285 ;
      RECT 164.595 21.24 165.7 21.41 ;
      RECT 164.83 19.655 165.395 20.625 ;
      RECT 164.935 18.415 165.395 20.625 ;
      RECT 164.83 18.415 165.395 18.985 ;
      RECT 164.475 22.645 165 22.865 ;
      RECT 164.83 21.58 165 22.865 ;
      RECT 164.83 21.58 165.36 21.945 ;
      RECT 163.875 19.945 164.135 20.625 ;
      RECT 163.875 19.945 164.66 20.165 ;
      RECT 164.46 18.875 164.66 20.165 ;
      RECT 164.46 19.155 164.765 19.485 ;
      RECT 163.875 18.875 164.66 19.045 ;
      RECT 163.875 18.415 164.135 19.045 ;
      RECT 164.135 23.065 164.47 23.235 ;
      RECT 164.135 22.795 164.305 23.235 ;
      RECT 164.08 21.56 164.25 22.925 ;
      RECT 164.135 21.135 164.385 21.69 ;
      RECT 163.415 20.295 163.685 20.625 ;
      RECT 163.515 18.415 163.685 20.625 ;
      RECT 163.515 19.215 164.29 19.775 ;
      RECT 163.415 18.415 163.685 18.745 ;
      RECT 162.345 19.945 162.745 20.625 ;
      RECT 162.345 19.945 163.29 20.165 ;
      RECT 163.055 18.875 163.29 20.165 ;
      RECT 163.055 19.155 163.345 19.485 ;
      RECT 162.345 18.875 163.29 19.045 ;
      RECT 162.345 18.415 162.745 19.045 ;
      RECT 162.435 22.795 162.605 23.255 ;
      RECT 162.435 22.795 163.1 22.965 ;
      RECT 162.87 21.635 163.1 22.965 ;
      RECT 162.435 21.635 163.1 21.805 ;
      RECT 162.435 21.135 162.605 21.805 ;
      RECT 160.415 17.335 160.745 17.855 ;
      RECT 160.625 16.585 160.795 17.42 ;
      RECT 160.57 17.295 160.795 17.42 ;
      RECT 160.58 16.585 160.795 16.715 ;
      RECT 160.405 15.74 160.735 16.665 ;
      RECT 160.415 22.775 160.745 23.295 ;
      RECT 160.625 22.025 160.795 22.86 ;
      RECT 160.57 22.735 160.795 22.86 ;
      RECT 160.58 22.025 160.795 22.155 ;
      RECT 160.405 21.18 160.735 22.105 ;
      RECT 159.575 17.335 159.905 17.86 ;
      RECT 159.705 16.835 159.905 17.86 ;
      RECT 159.705 16.835 160.455 17.165 ;
      RECT 159.705 15.695 159.895 17.86 ;
      RECT 159 16.255 159.895 16.63 ;
      RECT 159.555 15.695 159.895 16.63 ;
      RECT 159.575 22.775 159.905 23.3 ;
      RECT 159.705 22.275 159.905 23.3 ;
      RECT 159.705 22.275 160.455 22.605 ;
      RECT 159.705 21.135 159.895 23.3 ;
      RECT 159 21.695 159.895 22.07 ;
      RECT 159.555 21.135 159.895 22.07 ;
      RECT 159.945 19.655 160.275 20.58 ;
      RECT 160.165 18.9 160.335 19.735 ;
      RECT 160.12 19.605 160.335 19.735 ;
      RECT 160.11 18.9 160.335 19.025 ;
      RECT 159.955 18.465 160.285 18.985 ;
      RECT 160.06 28.455 160.315 28.785 ;
      RECT 160.145 26.575 160.315 28.785 ;
      RECT 160.13 28.375 160.315 28.785 ;
      RECT 160.06 26.575 160.315 27.245 ;
      RECT 159.095 19.69 159.435 20.625 ;
      RECT 159.245 18.46 159.435 20.625 ;
      RECT 158.54 19.69 159.435 20.065 ;
      RECT 159.245 19.155 159.995 19.485 ;
      RECT 159.245 18.46 159.445 19.485 ;
      RECT 159.115 18.46 159.445 18.985 ;
      RECT 157.81 28.535 159.345 28.785 ;
      RECT 159.175 28.135 159.345 28.785 ;
      RECT 156.915 28.135 157.085 28.785 ;
      RECT 157.81 28.135 157.98 28.785 ;
      RECT 159.175 28.135 159.975 28.305 ;
      RECT 159.805 27.415 159.975 28.305 ;
      RECT 156.915 28.135 157.98 28.305 ;
      RECT 156.915 27.415 159.975 27.585 ;
      RECT 156.915 26.575 157.085 27.585 ;
      RECT 159.21 27.765 159.575 27.965 ;
      RECT 159.21 27.765 159.585 27.935 ;
      RECT 158.045 17.625 158.83 17.795 ;
      RECT 158.66 15.825 158.83 17.795 ;
      RECT 158.66 16.835 159.535 17.165 ;
      RECT 157.945 15.825 158.83 15.995 ;
      RECT 158.045 23.065 158.83 23.235 ;
      RECT 158.66 21.265 158.83 23.235 ;
      RECT 158.66 22.275 159.535 22.605 ;
      RECT 157.945 21.265 158.83 21.435 ;
      RECT 157.755 27.005 159.39 27.245 ;
      RECT 159.14 26.575 159.39 27.245 ;
      RECT 157.755 26.915 157.985 27.245 ;
      RECT 157.485 20.325 158.37 20.495 ;
      RECT 158.2 18.525 158.37 20.495 ;
      RECT 158.2 19.155 159.075 19.485 ;
      RECT 157.585 18.525 158.37 18.695 ;
      RECT 158.71 27.765 158.995 28.365 ;
      RECT 158.71 27.765 159.04 27.965 ;
      RECT 158.025 17.125 158.49 17.455 ;
      RECT 158.17 16.165 158.49 17.455 ;
      RECT 158.025 22.565 158.49 22.895 ;
      RECT 158.17 21.605 158.49 22.895 ;
      RECT 158.16 27.765 158.44 28.365 ;
      RECT 157.965 27.765 158.44 27.965 ;
      RECT 157.255 26.575 157.585 27.245 ;
      RECT 158.095 26.575 158.425 26.785 ;
      RECT 157.255 26.575 158.425 26.745 ;
      RECT 158.235 25.055 158.405 26.065 ;
      RECT 155.345 25.055 158.405 25.225 ;
      RECT 155.345 24.335 155.515 25.225 ;
      RECT 157.34 24.335 158.405 24.505 ;
      RECT 158.235 23.855 158.405 24.505 ;
      RECT 155.345 24.335 156.145 24.505 ;
      RECT 155.975 23.855 156.145 24.505 ;
      RECT 157.34 23.855 157.51 24.505 ;
      RECT 155.975 23.855 157.51 24.105 ;
      RECT 156.895 25.895 158.065 26.065 ;
      RECT 157.735 25.395 158.065 26.065 ;
      RECT 156.895 25.855 157.225 26.065 ;
      RECT 157.71 18.865 158.03 20.155 ;
      RECT 157.565 18.865 158.03 19.195 ;
      RECT 157.47 17.625 157.875 17.795 ;
      RECT 157.47 15.695 157.64 17.795 ;
      RECT 156.81 17.095 157.64 17.395 ;
      RECT 156.81 17.065 157.01 17.395 ;
      RECT 157.47 15.695 157.72 16.025 ;
      RECT 157.47 23.065 157.875 23.235 ;
      RECT 157.47 21.135 157.64 23.235 ;
      RECT 156.81 22.535 157.64 22.835 ;
      RECT 156.81 22.505 157.01 22.835 ;
      RECT 157.47 21.135 157.72 21.465 ;
      RECT 155.93 25.395 156.18 26.065 ;
      RECT 157.335 25.395 157.565 25.725 ;
      RECT 155.93 25.395 157.565 25.635 ;
      RECT 157.01 20.295 157.26 20.625 ;
      RECT 157.01 18.525 157.18 20.625 ;
      RECT 156.35 18.925 156.55 19.255 ;
      RECT 156.35 18.925 157.18 19.225 ;
      RECT 157.01 18.525 157.415 18.695 ;
      RECT 156.88 24.675 157.355 24.875 ;
      RECT 156.88 24.275 157.16 24.875 ;
      RECT 155.925 17.625 156.6 17.795 ;
      RECT 156.43 16.675 156.6 17.795 ;
      RECT 157.13 16.585 157.3 16.915 ;
      RECT 156.43 16.675 157.3 16.845 ;
      RECT 156.79 16.585 157.3 16.845 ;
      RECT 156.79 15.8 156.96 16.845 ;
      RECT 155.855 15.8 156.96 15.97 ;
      RECT 155.925 23.065 156.6 23.235 ;
      RECT 156.43 22.115 156.6 23.235 ;
      RECT 157.13 22.025 157.3 22.355 ;
      RECT 156.43 22.115 157.3 22.285 ;
      RECT 156.79 22.025 157.3 22.285 ;
      RECT 156.79 21.24 156.96 22.285 ;
      RECT 155.855 21.24 156.96 21.41 ;
      RECT 155.395 20.35 156.5 20.52 ;
      RECT 156.33 19.475 156.5 20.52 ;
      RECT 156.33 19.475 156.84 19.735 ;
      RECT 156.67 19.405 156.84 19.735 ;
      RECT 155.97 19.475 156.84 19.645 ;
      RECT 155.97 18.525 156.14 19.645 ;
      RECT 155.465 18.525 156.14 18.695 ;
      RECT 155.735 17.205 156.26 17.425 ;
      RECT 156.09 16.14 156.26 17.425 ;
      RECT 156.09 16.14 156.62 16.505 ;
      RECT 155.735 22.645 156.26 22.865 ;
      RECT 156.09 21.58 156.26 22.865 ;
      RECT 156.09 21.58 156.62 21.945 ;
      RECT 156.28 24.675 156.61 24.875 ;
      RECT 156.325 24.275 156.61 24.875 ;
      RECT 155.63 19.815 156.16 20.18 ;
      RECT 155.63 18.895 155.8 20.18 ;
      RECT 155.275 18.895 155.8 19.115 ;
      RECT 155.735 24.705 156.11 24.875 ;
      RECT 155.745 24.675 156.11 24.875 ;
      RECT 155.395 17.625 155.73 17.795 ;
      RECT 155.395 17.355 155.565 17.795 ;
      RECT 155.34 16.12 155.51 17.485 ;
      RECT 155.395 15.695 155.645 16.25 ;
      RECT 155.395 23.065 155.73 23.235 ;
      RECT 155.395 22.795 155.565 23.235 ;
      RECT 155.34 21.56 155.51 22.925 ;
      RECT 155.395 21.135 155.645 21.69 ;
      RECT 154.935 20.07 155.185 20.625 ;
      RECT 154.88 18.835 155.05 20.2 ;
      RECT 154.935 18.525 155.105 18.965 ;
      RECT 154.935 18.525 155.27 18.695 ;
      RECT 155.005 25.395 155.26 26.065 ;
      RECT 155.005 23.855 155.175 26.065 ;
      RECT 155.005 23.855 155.19 24.265 ;
      RECT 155.005 23.855 155.215 24.195 ;
      RECT 155.005 23.855 155.26 24.185 ;
      RECT 153.695 17.355 153.865 17.815 ;
      RECT 153.695 17.355 154.36 17.525 ;
      RECT 154.13 16.195 154.36 17.525 ;
      RECT 153.695 16.195 154.36 16.365 ;
      RECT 153.695 15.695 153.865 16.365 ;
      RECT 153.695 22.795 153.865 23.255 ;
      RECT 153.695 22.795 154.36 22.965 ;
      RECT 154.13 21.635 154.36 22.965 ;
      RECT 153.695 21.635 154.36 21.805 ;
      RECT 153.695 21.135 153.865 21.805 ;
      RECT 153.235 19.955 153.405 20.625 ;
      RECT 153.235 19.955 153.9 20.125 ;
      RECT 153.67 18.795 153.9 20.125 ;
      RECT 153.235 18.795 153.9 18.965 ;
      RECT 153.235 18.505 153.405 18.965 ;
      RECT 152.635 25.045 152.965 26.065 ;
      RECT 151.795 25.045 152.125 26.065 ;
      RECT 151.465 25.045 152.965 25.215 ;
      RECT 151.465 24.335 151.64 25.215 ;
      RECT 149.015 24.675 151.64 24.845 ;
      RECT 151.465 24.335 152.885 24.505 ;
      RECT 152.715 23.855 152.885 24.505 ;
      RECT 151.875 23.86 152.045 24.505 ;
      RECT 148.635 11.815 148.805 12.465 ;
      RECT 149.475 11.815 149.645 12.46 ;
      RECT 148.635 11.815 150.055 11.985 ;
      RECT 149.88 11.105 150.055 11.985 ;
      RECT 149.88 11.475 152.505 11.645 ;
      RECT 148.555 11.105 150.055 11.275 ;
      RECT 149.395 10.255 149.725 11.275 ;
      RECT 148.555 10.255 148.885 11.275 ;
      RECT 145.8 17.575 146.055 17.905 ;
      RECT 145.885 15.695 146.055 17.905 ;
      RECT 145.845 17.565 146.055 17.905 ;
      RECT 145.87 17.495 146.055 17.905 ;
      RECT 145.8 15.695 146.055 16.365 ;
      RECT 145.8 19.955 146.055 20.625 ;
      RECT 145.885 18.415 146.055 20.625 ;
      RECT 145.87 18.415 146.055 18.825 ;
      RECT 145.845 18.415 146.055 18.755 ;
      RECT 145.8 18.415 146.055 18.745 ;
      RECT 143.55 17.655 145.085 17.905 ;
      RECT 144.915 17.255 145.085 17.905 ;
      RECT 142.655 17.255 142.825 17.905 ;
      RECT 143.55 17.255 143.72 17.905 ;
      RECT 144.915 17.255 145.715 17.425 ;
      RECT 145.545 16.535 145.715 17.425 ;
      RECT 142.655 17.255 143.72 17.425 ;
      RECT 142.655 16.535 145.715 16.705 ;
      RECT 142.655 15.695 142.825 16.705 ;
      RECT 142.655 19.615 142.825 20.625 ;
      RECT 142.655 19.615 145.715 19.785 ;
      RECT 145.545 18.895 145.715 19.785 ;
      RECT 144.915 18.895 145.715 19.065 ;
      RECT 142.655 18.895 143.72 19.065 ;
      RECT 143.55 18.415 143.72 19.065 ;
      RECT 144.915 18.415 145.085 19.065 ;
      RECT 142.655 18.415 142.825 19.065 ;
      RECT 143.55 18.415 145.085 18.665 ;
      RECT 144.95 16.885 145.315 17.085 ;
      RECT 144.95 16.885 145.375 17.055 ;
      RECT 144.95 19.265 145.325 19.435 ;
      RECT 144.95 19.235 145.315 19.435 ;
      RECT 143.495 16.125 145.13 16.365 ;
      RECT 144.88 15.695 145.13 16.365 ;
      RECT 143.495 16.035 143.725 16.365 ;
      RECT 144.88 19.955 145.13 20.625 ;
      RECT 143.495 19.955 143.725 20.285 ;
      RECT 143.495 19.955 145.13 20.195 ;
      RECT 144.45 16.885 144.735 17.485 ;
      RECT 144.45 16.885 144.78 17.085 ;
      RECT 144.45 19.235 144.78 19.435 ;
      RECT 144.45 18.835 144.735 19.435 ;
      RECT 144.355 14.165 144.685 15.185 ;
      RECT 143.515 14.165 143.845 15.185 ;
      RECT 143.185 14.165 144.685 14.335 ;
      RECT 143.185 13.455 143.36 14.335 ;
      RECT 140.735 13.795 143.36 13.965 ;
      RECT 143.185 13.455 144.605 13.625 ;
      RECT 144.435 12.975 144.605 13.625 ;
      RECT 143.595 12.98 143.765 13.625 ;
      RECT 143.9 16.885 144.18 17.485 ;
      RECT 143.705 16.885 144.18 17.085 ;
      RECT 143.705 19.235 144.18 19.435 ;
      RECT 143.9 18.835 144.18 19.435 ;
      RECT 142.995 15.695 143.325 16.365 ;
      RECT 143.835 15.695 144.165 15.905 ;
      RECT 142.995 15.695 144.165 15.865 ;
      RECT 142.995 20.455 144.165 20.625 ;
      RECT 143.835 20.415 144.165 20.625 ;
      RECT 142.995 19.955 143.325 20.625 ;
      RECT 142.015 28.215 142.345 28.735 ;
      RECT 142.225 27.465 142.395 28.3 ;
      RECT 142.17 28.175 142.395 28.3 ;
      RECT 142.18 27.465 142.395 27.595 ;
      RECT 142.005 26.62 142.335 27.545 ;
      RECT 138.515 11.815 138.685 12.465 ;
      RECT 139.355 11.815 139.525 12.46 ;
      RECT 138.515 11.815 139.935 11.985 ;
      RECT 139.76 11.105 139.935 11.985 ;
      RECT 139.76 11.475 142.385 11.645 ;
      RECT 138.435 11.105 139.935 11.275 ;
      RECT 139.275 10.255 139.605 11.275 ;
      RECT 138.435 10.255 138.765 11.275 ;
      RECT 141.175 28.215 141.505 28.74 ;
      RECT 141.305 27.715 141.505 28.74 ;
      RECT 141.305 27.715 142.055 28.045 ;
      RECT 141.305 26.575 141.495 28.74 ;
      RECT 140.6 27.135 141.495 27.51 ;
      RECT 141.155 26.575 141.495 27.51 ;
      RECT 141.555 22.775 141.885 23.295 ;
      RECT 141.765 22.025 141.935 22.86 ;
      RECT 141.71 22.735 141.935 22.86 ;
      RECT 141.72 22.025 141.935 22.155 ;
      RECT 141.545 21.18 141.875 22.105 ;
      RECT 140.715 22.775 141.045 23.3 ;
      RECT 140.845 22.275 141.045 23.3 ;
      RECT 140.845 22.275 141.595 22.605 ;
      RECT 140.845 21.135 141.035 23.3 ;
      RECT 140.14 21.695 141.035 22.07 ;
      RECT 140.695 21.135 141.035 22.07 ;
      RECT 141.215 25.055 141.385 26.065 ;
      RECT 138.325 25.055 141.385 25.225 ;
      RECT 138.325 24.335 138.495 25.225 ;
      RECT 140.32 24.335 141.385 24.505 ;
      RECT 141.215 23.855 141.385 24.505 ;
      RECT 138.325 24.335 139.125 24.505 ;
      RECT 138.955 23.855 139.125 24.505 ;
      RECT 140.32 23.855 140.49 24.505 ;
      RECT 138.955 23.855 140.49 24.105 ;
      RECT 141.215 30.495 141.385 31.505 ;
      RECT 138.325 30.495 141.385 30.665 ;
      RECT 138.325 29.775 138.495 30.665 ;
      RECT 140.32 29.775 141.385 29.945 ;
      RECT 141.215 29.295 141.385 29.945 ;
      RECT 138.325 29.775 139.125 29.945 ;
      RECT 138.955 29.295 139.125 29.945 ;
      RECT 140.32 29.295 140.49 29.945 ;
      RECT 138.955 29.295 140.49 29.545 ;
      RECT 139.645 28.505 140.43 28.675 ;
      RECT 140.26 26.705 140.43 28.675 ;
      RECT 140.26 27.715 141.135 28.045 ;
      RECT 139.545 26.705 140.43 26.875 ;
      RECT 139.875 25.895 141.045 26.065 ;
      RECT 140.715 25.395 141.045 26.065 ;
      RECT 139.875 25.855 140.205 26.065 ;
      RECT 139.875 31.335 141.045 31.505 ;
      RECT 140.715 30.835 141.045 31.505 ;
      RECT 139.875 31.295 140.205 31.505 ;
      RECT 139.185 23.065 139.97 23.235 ;
      RECT 139.8 21.265 139.97 23.235 ;
      RECT 139.8 22.275 140.675 22.605 ;
      RECT 139.085 21.265 139.97 21.435 ;
      RECT 138.91 25.395 139.16 26.065 ;
      RECT 140.315 25.395 140.545 25.725 ;
      RECT 138.91 25.395 140.545 25.635 ;
      RECT 138.91 30.835 139.16 31.505 ;
      RECT 140.315 30.835 140.545 31.165 ;
      RECT 138.91 30.835 140.545 31.075 ;
      RECT 139.86 24.675 140.335 24.875 ;
      RECT 139.86 24.275 140.14 24.875 ;
      RECT 139.86 30.115 140.335 30.315 ;
      RECT 139.86 29.715 140.14 30.315 ;
      RECT 139.705 19.655 140.035 20.58 ;
      RECT 139.925 18.9 140.095 19.735 ;
      RECT 139.88 19.605 140.095 19.735 ;
      RECT 139.87 18.9 140.095 19.025 ;
      RECT 139.715 18.465 140.045 18.985 ;
      RECT 139.625 28.005 140.09 28.335 ;
      RECT 139.77 27.045 140.09 28.335 ;
      RECT 138.855 19.69 139.195 20.625 ;
      RECT 139.005 18.46 139.195 20.625 ;
      RECT 138.3 19.69 139.195 20.065 ;
      RECT 139.005 19.155 139.755 19.485 ;
      RECT 139.005 18.46 139.205 19.485 ;
      RECT 138.875 18.46 139.205 18.985 ;
      RECT 139.165 22.565 139.63 22.895 ;
      RECT 139.31 21.605 139.63 22.895 ;
      RECT 139.26 24.675 139.59 24.875 ;
      RECT 139.305 24.275 139.59 24.875 ;
      RECT 139.26 30.115 139.59 30.315 ;
      RECT 139.305 29.715 139.59 30.315 ;
      RECT 139.07 28.505 139.475 28.675 ;
      RECT 139.07 26.575 139.24 28.675 ;
      RECT 138.41 27.975 139.24 28.275 ;
      RECT 138.41 27.945 138.61 28.275 ;
      RECT 139.07 26.575 139.32 26.905 ;
      RECT 138.715 24.705 139.09 24.875 ;
      RECT 138.725 24.675 139.09 24.875 ;
      RECT 138.715 30.145 139.09 30.315 ;
      RECT 138.725 30.115 139.09 30.315 ;
      RECT 138.61 23.065 139.015 23.235 ;
      RECT 138.61 21.135 138.78 23.235 ;
      RECT 137.95 22.535 138.78 22.835 ;
      RECT 137.95 22.505 138.15 22.835 ;
      RECT 138.61 21.135 138.86 21.465 ;
      RECT 137.525 28.505 138.2 28.675 ;
      RECT 138.03 27.555 138.2 28.675 ;
      RECT 138.73 27.465 138.9 27.795 ;
      RECT 138.03 27.555 138.9 27.725 ;
      RECT 138.39 27.465 138.9 27.725 ;
      RECT 138.39 26.68 138.56 27.725 ;
      RECT 137.455 26.68 138.56 26.85 ;
      RECT 137.245 20.325 138.13 20.495 ;
      RECT 137.96 18.525 138.13 20.495 ;
      RECT 137.96 19.155 138.835 19.485 ;
      RECT 137.345 18.525 138.13 18.695 ;
      RECT 137.065 23.065 137.74 23.235 ;
      RECT 137.57 22.115 137.74 23.235 ;
      RECT 138.27 22.025 138.44 22.355 ;
      RECT 137.57 22.115 138.44 22.285 ;
      RECT 137.93 22.025 138.44 22.285 ;
      RECT 137.93 21.24 138.1 22.285 ;
      RECT 136.995 21.24 138.1 21.41 ;
      RECT 137.985 25.395 138.24 26.065 ;
      RECT 137.985 23.855 138.155 26.065 ;
      RECT 137.985 23.855 138.17 24.265 ;
      RECT 137.985 23.855 138.195 24.195 ;
      RECT 137.985 23.855 138.24 24.185 ;
      RECT 137.985 30.835 138.24 31.505 ;
      RECT 137.985 29.295 138.155 31.505 ;
      RECT 137.985 29.295 138.17 29.705 ;
      RECT 137.985 29.295 138.195 29.635 ;
      RECT 137.985 29.295 138.24 29.625 ;
      RECT 137.98 17.575 138.235 17.905 ;
      RECT 138.065 15.695 138.235 17.905 ;
      RECT 138.025 17.565 138.235 17.905 ;
      RECT 138.05 17.495 138.235 17.905 ;
      RECT 137.98 15.695 138.235 16.365 ;
      RECT 137.335 28.085 137.86 28.305 ;
      RECT 137.69 27.02 137.86 28.305 ;
      RECT 137.69 27.02 138.22 27.385 ;
      RECT 135.73 17.655 137.265 17.905 ;
      RECT 137.095 17.255 137.265 17.905 ;
      RECT 134.835 17.255 135.005 17.905 ;
      RECT 135.73 17.255 135.9 17.905 ;
      RECT 137.095 17.255 137.895 17.425 ;
      RECT 137.725 16.535 137.895 17.425 ;
      RECT 134.835 17.255 135.9 17.425 ;
      RECT 134.835 16.535 137.895 16.705 ;
      RECT 134.835 15.695 135.005 16.705 ;
      RECT 137.47 18.865 137.79 20.155 ;
      RECT 137.325 18.865 137.79 19.195 ;
      RECT 136.875 22.645 137.4 22.865 ;
      RECT 137.23 21.58 137.4 22.865 ;
      RECT 137.23 21.58 137.76 21.945 ;
      RECT 137.13 16.885 137.495 17.085 ;
      RECT 137.13 16.885 137.505 17.055 ;
      RECT 136.995 28.505 137.33 28.675 ;
      RECT 136.995 28.235 137.165 28.675 ;
      RECT 136.94 27 137.11 28.365 ;
      RECT 136.995 26.575 137.245 27.13 ;
      RECT 135.675 16.125 137.31 16.365 ;
      RECT 137.06 15.695 137.31 16.365 ;
      RECT 135.675 16.035 135.905 16.365 ;
      RECT 136.77 20.295 137.02 20.625 ;
      RECT 136.77 18.525 136.94 20.625 ;
      RECT 136.11 18.925 136.31 19.255 ;
      RECT 136.11 18.925 136.94 19.225 ;
      RECT 136.77 18.525 137.175 18.695 ;
      RECT 136.63 16.885 136.915 17.485 ;
      RECT 136.63 16.885 136.96 17.085 ;
      RECT 136.57 16.885 136.96 17.055 ;
      RECT 136.535 23.065 136.87 23.235 ;
      RECT 136.535 22.795 136.705 23.235 ;
      RECT 136.48 21.56 136.65 22.925 ;
      RECT 136.535 21.135 136.785 21.69 ;
      RECT 133.755 14.165 134.085 15.185 ;
      RECT 132.915 14.165 133.245 15.185 ;
      RECT 132.915 14.165 134.415 14.335 ;
      RECT 134.24 13.455 134.415 14.335 ;
      RECT 134.24 13.795 136.865 13.965 ;
      RECT 132.995 13.455 134.415 13.625 ;
      RECT 133.835 12.98 134.005 13.625 ;
      RECT 132.995 12.975 133.165 13.625 ;
      RECT 135.155 20.35 136.26 20.52 ;
      RECT 136.09 19.475 136.26 20.52 ;
      RECT 136.09 19.475 136.6 19.735 ;
      RECT 136.43 19.405 136.6 19.735 ;
      RECT 135.73 19.475 136.6 19.645 ;
      RECT 135.73 18.525 135.9 19.645 ;
      RECT 135.225 18.525 135.9 18.695 ;
      RECT 136.08 16.885 136.36 17.485 ;
      RECT 135.885 16.885 136.36 17.085 ;
      RECT 135.175 15.695 135.505 16.365 ;
      RECT 136.015 15.695 136.345 15.905 ;
      RECT 135.175 15.695 136.345 15.865 ;
      RECT 135.295 28.235 135.465 28.695 ;
      RECT 135.295 28.235 135.96 28.405 ;
      RECT 135.73 27.075 135.96 28.405 ;
      RECT 135.295 27.075 135.96 27.245 ;
      RECT 135.295 26.575 135.465 27.245 ;
      RECT 135.39 19.815 135.92 20.18 ;
      RECT 135.39 18.895 135.56 20.18 ;
      RECT 135.035 18.895 135.56 19.115 ;
      RECT 134.835 22.795 135.005 23.255 ;
      RECT 134.835 22.795 135.5 22.965 ;
      RECT 135.27 21.635 135.5 22.965 ;
      RECT 134.835 21.635 135.5 21.805 ;
      RECT 134.835 21.135 135.005 21.805 ;
      RECT 134.695 20.07 134.945 20.625 ;
      RECT 134.64 18.835 134.81 20.2 ;
      RECT 134.695 18.525 134.865 18.965 ;
      RECT 134.695 18.525 135.03 18.695 ;
      RECT 134.315 22.84 134.575 23.345 ;
      RECT 134.405 21.135 134.575 23.345 ;
      RECT 134.305 21.135 134.575 22.04 ;
      RECT 133.455 22.795 133.625 23.345 ;
      RECT 133.455 22.795 134.12 22.965 ;
      RECT 133.95 21.895 134.12 22.965 ;
      RECT 133.95 22.21 134.235 22.54 ;
      RECT 133.455 21.895 134.12 22.065 ;
      RECT 133.455 21.135 133.625 22.065 ;
      RECT 132.995 19.955 133.165 20.625 ;
      RECT 132.995 19.955 133.66 20.125 ;
      RECT 133.43 18.795 133.66 20.125 ;
      RECT 132.995 18.795 133.66 18.965 ;
      RECT 132.995 18.505 133.165 18.965 ;
      RECT 131.435 22.775 131.765 23.295 ;
      RECT 131.645 22.025 131.815 22.86 ;
      RECT 131.59 22.735 131.815 22.86 ;
      RECT 131.6 22.025 131.815 22.155 ;
      RECT 131.425 21.18 131.755 22.105 ;
      RECT 131.435 28.215 131.765 28.735 ;
      RECT 131.645 27.465 131.815 28.3 ;
      RECT 131.59 28.175 131.815 28.3 ;
      RECT 131.6 27.465 131.815 27.595 ;
      RECT 131.425 26.62 131.755 27.545 ;
      RECT 130.595 22.775 130.925 23.3 ;
      RECT 130.725 22.275 130.925 23.3 ;
      RECT 130.725 22.275 131.475 22.605 ;
      RECT 130.725 21.135 130.915 23.3 ;
      RECT 130.02 21.695 130.915 22.07 ;
      RECT 130.575 21.135 130.915 22.07 ;
      RECT 130.595 28.215 130.925 28.74 ;
      RECT 130.725 27.715 130.925 28.74 ;
      RECT 130.725 27.715 131.475 28.045 ;
      RECT 130.725 26.575 130.915 28.74 ;
      RECT 130.02 27.135 130.915 27.51 ;
      RECT 130.575 26.575 130.915 27.51 ;
      RECT 129.065 23.065 129.85 23.235 ;
      RECT 129.68 21.265 129.85 23.235 ;
      RECT 129.68 22.275 130.555 22.605 ;
      RECT 128.965 21.265 129.85 21.435 ;
      RECT 129.065 28.505 129.85 28.675 ;
      RECT 129.68 26.705 129.85 28.675 ;
      RECT 129.68 27.715 130.555 28.045 ;
      RECT 128.965 26.705 129.85 26.875 ;
      RECT 129.045 22.565 129.51 22.895 ;
      RECT 129.19 21.605 129.51 22.895 ;
      RECT 129.045 28.005 129.51 28.335 ;
      RECT 129.19 27.045 129.51 28.335 ;
      RECT 128.78 17.575 129.035 17.905 ;
      RECT 128.865 15.695 129.035 17.905 ;
      RECT 128.825 17.565 129.035 17.905 ;
      RECT 128.85 17.495 129.035 17.905 ;
      RECT 128.78 15.695 129.035 16.365 ;
      RECT 128.49 23.065 128.895 23.235 ;
      RECT 128.49 21.135 128.66 23.235 ;
      RECT 127.83 22.535 128.66 22.835 ;
      RECT 127.83 22.505 128.03 22.835 ;
      RECT 128.49 21.135 128.74 21.465 ;
      RECT 128.49 28.505 128.895 28.675 ;
      RECT 128.49 26.575 128.66 28.675 ;
      RECT 127.83 27.975 128.66 28.275 ;
      RECT 127.83 27.945 128.03 28.275 ;
      RECT 128.49 26.575 128.74 26.905 ;
      RECT 126.53 17.655 128.065 17.905 ;
      RECT 127.895 17.255 128.065 17.905 ;
      RECT 125.635 17.255 125.805 17.905 ;
      RECT 126.53 17.255 126.7 17.905 ;
      RECT 127.895 17.255 128.695 17.425 ;
      RECT 128.525 16.535 128.695 17.425 ;
      RECT 125.635 17.255 126.7 17.425 ;
      RECT 125.635 16.535 128.695 16.705 ;
      RECT 125.635 15.695 125.805 16.705 ;
      RECT 126.945 23.065 127.62 23.235 ;
      RECT 127.45 22.115 127.62 23.235 ;
      RECT 128.15 22.025 128.32 22.355 ;
      RECT 127.45 22.115 128.32 22.285 ;
      RECT 127.81 22.025 128.32 22.285 ;
      RECT 127.81 21.24 127.98 22.285 ;
      RECT 126.875 21.24 127.98 21.41 ;
      RECT 126.945 28.505 127.62 28.675 ;
      RECT 127.45 27.555 127.62 28.675 ;
      RECT 128.15 27.465 128.32 27.795 ;
      RECT 127.45 27.555 128.32 27.725 ;
      RECT 127.81 27.465 128.32 27.725 ;
      RECT 127.81 26.68 127.98 27.725 ;
      RECT 126.875 26.68 127.98 26.85 ;
      RECT 127.93 16.885 128.295 17.085 ;
      RECT 127.93 16.885 128.305 17.055 ;
      RECT 126.475 16.125 128.11 16.365 ;
      RECT 127.86 15.695 128.11 16.365 ;
      RECT 126.475 16.035 126.705 16.365 ;
      RECT 127.43 16.885 127.715 17.485 ;
      RECT 127.43 16.885 127.76 17.085 ;
      RECT 126.755 22.645 127.28 22.865 ;
      RECT 127.11 21.58 127.28 22.865 ;
      RECT 127.11 21.58 127.64 21.945 ;
      RECT 126.755 28.085 127.28 28.305 ;
      RECT 127.11 27.02 127.28 28.305 ;
      RECT 127.11 27.02 127.64 27.385 ;
      RECT 126.88 16.885 127.16 17.485 ;
      RECT 126.685 16.885 127.16 17.085 ;
      RECT 125.975 15.695 126.305 16.365 ;
      RECT 126.815 15.695 127.145 15.905 ;
      RECT 125.975 15.695 127.145 15.865 ;
      RECT 126.415 23.065 126.75 23.235 ;
      RECT 126.415 22.795 126.585 23.235 ;
      RECT 126.36 21.56 126.53 22.925 ;
      RECT 126.415 21.135 126.665 21.69 ;
      RECT 126.415 28.505 126.75 28.675 ;
      RECT 126.415 28.235 126.585 28.675 ;
      RECT 126.36 27 126.53 28.365 ;
      RECT 126.415 26.575 126.665 27.13 ;
      RECT 124.715 22.795 124.885 23.255 ;
      RECT 124.715 22.795 125.38 22.965 ;
      RECT 125.15 21.635 125.38 22.965 ;
      RECT 124.715 21.635 125.38 21.805 ;
      RECT 124.715 21.135 124.885 21.805 ;
      RECT 124.715 28.235 124.885 28.695 ;
      RECT 124.715 28.235 125.38 28.405 ;
      RECT 125.15 27.075 125.38 28.405 ;
      RECT 124.715 27.075 125.38 27.245 ;
      RECT 124.715 26.575 124.885 27.245 ;
      RECT 124.985 19.655 125.315 20.58 ;
      RECT 125.205 18.9 125.375 19.735 ;
      RECT 125.16 19.605 125.375 19.735 ;
      RECT 125.15 18.9 125.375 19.025 ;
      RECT 124.995 18.465 125.325 18.985 ;
      RECT 124.985 25.095 125.315 26.02 ;
      RECT 125.205 24.34 125.375 25.175 ;
      RECT 125.16 25.045 125.375 25.175 ;
      RECT 125.15 24.34 125.375 24.465 ;
      RECT 124.995 23.905 125.325 24.425 ;
      RECT 124.135 19.69 124.475 20.625 ;
      RECT 124.285 18.46 124.475 20.625 ;
      RECT 123.58 19.69 124.475 20.065 ;
      RECT 124.285 19.155 125.035 19.485 ;
      RECT 124.285 18.46 124.485 19.485 ;
      RECT 124.155 18.46 124.485 18.985 ;
      RECT 124.135 25.13 124.475 26.065 ;
      RECT 124.285 23.9 124.475 26.065 ;
      RECT 123.58 25.13 124.475 25.505 ;
      RECT 124.285 24.595 125.035 24.925 ;
      RECT 124.285 23.9 124.485 24.925 ;
      RECT 124.155 23.9 124.485 24.425 ;
      RECT 122.525 20.325 123.41 20.495 ;
      RECT 123.24 18.525 123.41 20.495 ;
      RECT 123.24 19.155 124.115 19.485 ;
      RECT 122.625 18.525 123.41 18.695 ;
      RECT 122.525 25.765 123.41 25.935 ;
      RECT 123.24 23.965 123.41 25.935 ;
      RECT 123.24 24.595 124.115 24.925 ;
      RECT 122.625 23.965 123.41 24.135 ;
      RECT 123.275 11.815 123.445 12.465 ;
      RECT 122.435 11.815 122.605 12.46 ;
      RECT 122.025 11.815 123.445 11.985 ;
      RECT 122.025 11.105 122.2 11.985 ;
      RECT 119.575 11.475 122.2 11.645 ;
      RECT 122.025 11.105 123.525 11.275 ;
      RECT 123.195 10.255 123.525 11.275 ;
      RECT 122.355 10.255 122.685 11.275 ;
      RECT 123.275 17.255 123.445 17.905 ;
      RECT 122.435 17.255 122.605 17.9 ;
      RECT 122.025 17.255 123.445 17.425 ;
      RECT 122.025 16.545 122.2 17.425 ;
      RECT 119.575 16.915 122.2 17.085 ;
      RECT 122.025 16.545 123.525 16.715 ;
      RECT 123.195 15.695 123.525 16.715 ;
      RECT 122.355 15.695 122.685 16.715 ;
      RECT 122.75 18.865 123.07 20.155 ;
      RECT 122.605 18.865 123.07 19.195 ;
      RECT 122.75 24.305 123.07 25.595 ;
      RECT 122.605 24.305 123.07 24.635 ;
      RECT 122.8 28.455 123.055 28.785 ;
      RECT 122.885 26.575 123.055 28.785 ;
      RECT 122.845 28.445 123.055 28.785 ;
      RECT 122.87 28.375 123.055 28.785 ;
      RECT 122.8 26.575 123.055 27.245 ;
      RECT 122.8 30.835 123.055 31.505 ;
      RECT 122.885 29.295 123.055 31.505 ;
      RECT 122.87 29.295 123.055 29.705 ;
      RECT 122.845 29.295 123.055 29.635 ;
      RECT 122.8 29.295 123.055 29.625 ;
      RECT 120.55 28.535 122.085 28.785 ;
      RECT 121.915 28.135 122.085 28.785 ;
      RECT 119.655 28.135 119.825 28.785 ;
      RECT 120.55 28.135 120.72 28.785 ;
      RECT 121.915 28.135 122.715 28.305 ;
      RECT 122.545 27.415 122.715 28.305 ;
      RECT 119.655 28.135 120.72 28.305 ;
      RECT 119.655 27.415 122.715 27.585 ;
      RECT 119.655 26.575 119.825 27.585 ;
      RECT 119.655 30.495 119.825 31.505 ;
      RECT 119.655 30.495 122.715 30.665 ;
      RECT 122.545 29.775 122.715 30.665 ;
      RECT 121.915 29.775 122.715 29.945 ;
      RECT 119.655 29.775 120.72 29.945 ;
      RECT 120.55 29.295 120.72 29.945 ;
      RECT 121.915 29.295 122.085 29.945 ;
      RECT 119.655 29.295 119.825 29.945 ;
      RECT 120.55 29.295 122.085 29.545 ;
      RECT 122.05 20.295 122.3 20.625 ;
      RECT 122.05 18.525 122.22 20.625 ;
      RECT 121.39 18.925 121.59 19.255 ;
      RECT 121.39 18.925 122.22 19.225 ;
      RECT 122.05 18.525 122.455 18.695 ;
      RECT 122.05 25.735 122.3 26.065 ;
      RECT 122.05 23.965 122.22 26.065 ;
      RECT 121.39 24.365 121.59 24.695 ;
      RECT 121.39 24.365 122.22 24.665 ;
      RECT 122.05 23.965 122.455 24.135 ;
      RECT 121.95 27.765 122.315 27.965 ;
      RECT 121.95 27.765 122.325 27.935 ;
      RECT 121.95 30.145 122.325 30.315 ;
      RECT 121.95 30.115 122.315 30.315 ;
      RECT 120.495 27.005 122.13 27.245 ;
      RECT 121.88 26.575 122.13 27.245 ;
      RECT 120.495 26.915 120.725 27.245 ;
      RECT 121.88 30.835 122.13 31.505 ;
      RECT 120.495 30.835 120.725 31.165 ;
      RECT 120.495 30.835 122.13 31.075 ;
      RECT 120.435 20.35 121.54 20.52 ;
      RECT 121.37 19.475 121.54 20.52 ;
      RECT 121.37 19.475 121.88 19.735 ;
      RECT 121.71 19.405 121.88 19.735 ;
      RECT 121.01 19.475 121.88 19.645 ;
      RECT 121.01 18.525 121.18 19.645 ;
      RECT 120.505 18.525 121.18 18.695 ;
      RECT 120.435 25.79 121.54 25.96 ;
      RECT 121.37 24.915 121.54 25.96 ;
      RECT 121.37 24.915 121.88 25.175 ;
      RECT 121.71 24.845 121.88 25.175 ;
      RECT 121.01 24.915 121.88 25.085 ;
      RECT 121.01 23.965 121.18 25.085 ;
      RECT 120.505 23.965 121.18 24.135 ;
      RECT 121.45 27.765 121.735 28.365 ;
      RECT 121.45 27.765 121.78 27.965 ;
      RECT 121.45 30.115 121.78 30.315 ;
      RECT 121.45 29.715 121.735 30.315 ;
      RECT 121.42 14.515 121.675 15.185 ;
      RECT 121.505 12.975 121.675 15.185 ;
      RECT 121.49 12.975 121.675 13.385 ;
      RECT 121.465 12.975 121.675 13.315 ;
      RECT 121.42 12.975 121.675 13.305 ;
      RECT 118.275 14.175 118.445 15.185 ;
      RECT 118.275 14.175 121.335 14.345 ;
      RECT 121.165 13.455 121.335 14.345 ;
      RECT 120.535 13.455 121.335 13.625 ;
      RECT 118.275 13.455 119.34 13.625 ;
      RECT 119.17 12.975 119.34 13.625 ;
      RECT 120.535 12.975 120.705 13.625 ;
      RECT 118.275 12.975 118.445 13.625 ;
      RECT 119.17 12.975 120.705 13.225 ;
      RECT 120.67 19.815 121.2 20.18 ;
      RECT 120.67 18.895 120.84 20.18 ;
      RECT 120.315 18.895 120.84 19.115 ;
      RECT 120.67 25.255 121.2 25.62 ;
      RECT 120.67 24.335 120.84 25.62 ;
      RECT 120.315 24.335 120.84 24.555 ;
      RECT 120.9 27.765 121.18 28.365 ;
      RECT 120.705 27.765 121.18 27.965 ;
      RECT 120.705 30.115 121.18 30.315 ;
      RECT 120.9 29.715 121.18 30.315 ;
      RECT 119.995 26.575 120.325 27.245 ;
      RECT 120.835 26.575 121.165 26.785 ;
      RECT 119.995 26.575 121.165 26.745 ;
      RECT 119.995 31.335 121.165 31.505 ;
      RECT 120.835 31.295 121.165 31.505 ;
      RECT 119.995 30.835 120.325 31.505 ;
      RECT 120.57 13.825 120.995 13.995 ;
      RECT 120.57 13.795 120.935 13.995 ;
      RECT 120.5 14.515 120.75 15.185 ;
      RECT 119.115 14.515 119.345 14.845 ;
      RECT 119.115 14.515 120.75 14.755 ;
      RECT 120.07 13.795 120.4 13.995 ;
      RECT 120.07 13.395 120.355 13.995 ;
      RECT 119.975 20.07 120.225 20.625 ;
      RECT 119.92 18.835 120.09 20.2 ;
      RECT 119.975 18.525 120.145 18.965 ;
      RECT 119.975 18.525 120.31 18.695 ;
      RECT 119.975 25.51 120.225 26.065 ;
      RECT 119.92 24.275 120.09 25.64 ;
      RECT 119.975 23.965 120.145 24.405 ;
      RECT 119.975 23.965 120.31 24.135 ;
      RECT 119.545 33.595 119.875 34.225 ;
      RECT 119.545 32.015 119.795 34.225 ;
      RECT 119.545 32.015 119.875 32.995 ;
      RECT 119.325 13.795 119.8 13.995 ;
      RECT 119.52 13.395 119.8 13.995 ;
      RECT 118.615 15.015 119.785 15.185 ;
      RECT 119.455 14.975 119.785 15.185 ;
      RECT 118.615 14.515 118.945 15.185 ;
      RECT 118.275 19.955 118.445 20.625 ;
      RECT 118.275 19.955 118.94 20.125 ;
      RECT 118.71 18.795 118.94 20.125 ;
      RECT 118.275 18.795 118.94 18.965 ;
      RECT 118.275 18.505 118.445 18.965 ;
      RECT 118.275 25.395 118.445 26.065 ;
      RECT 118.275 25.395 118.94 25.565 ;
      RECT 118.71 24.235 118.94 25.565 ;
      RECT 118.275 24.235 118.94 24.405 ;
      RECT 118.275 23.945 118.445 24.405 ;
      RECT 117.175 22.775 117.505 23.295 ;
      RECT 117.385 22.025 117.555 22.86 ;
      RECT 117.33 22.735 117.555 22.86 ;
      RECT 117.34 22.025 117.555 22.155 ;
      RECT 117.165 21.18 117.495 22.105 ;
      RECT 116.335 22.775 116.665 23.3 ;
      RECT 116.465 22.275 116.665 23.3 ;
      RECT 116.465 22.275 117.215 22.605 ;
      RECT 116.465 21.135 116.655 23.3 ;
      RECT 115.76 21.695 116.655 22.07 ;
      RECT 116.315 21.135 116.655 22.07 ;
      RECT 114.805 23.065 115.59 23.235 ;
      RECT 115.42 21.265 115.59 23.235 ;
      RECT 115.42 22.275 116.295 22.605 ;
      RECT 114.705 21.265 115.59 21.435 ;
      RECT 115.9 25.395 116.155 26.065 ;
      RECT 115.985 23.855 116.155 26.065 ;
      RECT 115.97 23.855 116.155 24.265 ;
      RECT 115.945 23.855 116.155 24.195 ;
      RECT 115.9 23.855 116.155 24.185 ;
      RECT 112.755 25.055 112.925 26.065 ;
      RECT 112.755 25.055 115.815 25.225 ;
      RECT 115.645 24.335 115.815 25.225 ;
      RECT 115.015 24.335 115.815 24.505 ;
      RECT 112.755 24.335 113.82 24.505 ;
      RECT 113.65 23.855 113.82 24.505 ;
      RECT 115.015 23.855 115.185 24.505 ;
      RECT 112.755 23.855 112.925 24.505 ;
      RECT 113.65 23.855 115.185 24.105 ;
      RECT 115.375 14.165 115.705 15.185 ;
      RECT 114.535 14.165 114.865 15.185 ;
      RECT 114.205 14.165 115.705 14.335 ;
      RECT 114.205 13.455 114.38 14.335 ;
      RECT 111.755 13.795 114.38 13.965 ;
      RECT 114.205 13.455 115.625 13.625 ;
      RECT 115.455 12.975 115.625 13.625 ;
      RECT 114.615 12.98 114.785 13.625 ;
      RECT 115.05 24.705 115.425 24.875 ;
      RECT 115.05 24.675 115.415 24.875 ;
      RECT 114.785 22.565 115.25 22.895 ;
      RECT 114.93 21.605 115.25 22.895 ;
      RECT 114.98 25.395 115.23 26.065 ;
      RECT 113.595 25.395 113.825 25.725 ;
      RECT 113.595 25.395 115.23 25.635 ;
      RECT 114.55 24.675 114.88 24.875 ;
      RECT 114.55 24.275 114.835 24.875 ;
      RECT 114.455 19.605 114.785 20.625 ;
      RECT 113.615 19.605 113.945 20.625 ;
      RECT 113.285 19.605 114.785 19.775 ;
      RECT 113.285 18.895 113.46 19.775 ;
      RECT 110.835 19.235 113.46 19.405 ;
      RECT 113.285 18.895 114.705 19.065 ;
      RECT 114.535 18.415 114.705 19.065 ;
      RECT 113.695 18.42 113.865 19.065 ;
      RECT 114.52 17.575 114.775 17.905 ;
      RECT 114.605 15.695 114.775 17.905 ;
      RECT 114.565 17.565 114.775 17.905 ;
      RECT 114.59 17.495 114.775 17.905 ;
      RECT 114.52 15.695 114.775 16.365 ;
      RECT 114.23 23.065 114.635 23.235 ;
      RECT 114.23 21.135 114.4 23.235 ;
      RECT 113.57 22.535 114.4 22.835 ;
      RECT 113.57 22.505 113.77 22.835 ;
      RECT 114.23 21.135 114.48 21.465 ;
      RECT 112.27 17.655 113.805 17.905 ;
      RECT 113.635 17.255 113.805 17.905 ;
      RECT 111.375 17.255 111.545 17.905 ;
      RECT 112.27 17.255 112.44 17.905 ;
      RECT 113.635 17.255 114.435 17.425 ;
      RECT 114.265 16.535 114.435 17.425 ;
      RECT 111.375 17.255 112.44 17.425 ;
      RECT 111.375 16.535 114.435 16.705 ;
      RECT 111.375 15.695 111.545 16.705 ;
      RECT 113.805 24.675 114.28 24.875 ;
      RECT 114 24.275 114.28 24.875 ;
      RECT 113.095 25.895 114.265 26.065 ;
      RECT 113.935 25.855 114.265 26.065 ;
      RECT 113.095 25.395 113.425 26.065 ;
      RECT 112.685 23.065 113.36 23.235 ;
      RECT 113.19 22.115 113.36 23.235 ;
      RECT 113.89 22.025 114.06 22.355 ;
      RECT 113.19 22.115 114.06 22.285 ;
      RECT 113.55 22.025 114.06 22.285 ;
      RECT 113.55 21.24 113.72 22.285 ;
      RECT 112.615 21.24 113.72 21.41 ;
      RECT 113.67 16.885 114.035 17.085 ;
      RECT 113.67 16.885 114.045 17.055 ;
      RECT 112.215 16.125 113.85 16.365 ;
      RECT 113.6 15.695 113.85 16.365 ;
      RECT 112.215 16.035 112.445 16.365 ;
      RECT 113.17 16.885 113.455 17.485 ;
      RECT 113.17 16.885 113.5 17.085 ;
      RECT 112.495 22.645 113.02 22.865 ;
      RECT 112.85 21.58 113.02 22.865 ;
      RECT 112.85 21.58 113.38 21.945 ;
      RECT 112.62 16.885 112.9 17.485 ;
      RECT 112.425 16.885 112.9 17.085 ;
      RECT 111.715 15.695 112.045 16.365 ;
      RECT 112.555 15.695 112.885 15.905 ;
      RECT 111.715 15.695 112.885 15.865 ;
      RECT 112.155 23.065 112.49 23.235 ;
      RECT 112.155 22.795 112.325 23.235 ;
      RECT 112.1 21.56 112.27 22.925 ;
      RECT 112.155 21.135 112.405 21.69 ;
      RECT 110.455 22.795 110.625 23.255 ;
      RECT 110.455 22.795 111.12 22.965 ;
      RECT 110.89 21.635 111.12 22.965 ;
      RECT 110.455 21.635 111.12 21.805 ;
      RECT 110.455 21.135 110.625 21.805 ;
      RECT 104.315 14.165 104.645 15.185 ;
      RECT 103.475 14.165 103.805 15.185 ;
      RECT 103.475 14.165 104.975 14.335 ;
      RECT 104.8 13.455 104.975 14.335 ;
      RECT 104.8 13.795 107.425 13.965 ;
      RECT 103.555 13.455 104.975 13.625 ;
      RECT 104.395 12.98 104.565 13.625 ;
      RECT 103.555 12.975 103.725 13.625 ;
      RECT 103.555 17.255 103.725 17.905 ;
      RECT 104.395 17.255 104.565 17.9 ;
      RECT 103.555 17.255 104.975 17.425 ;
      RECT 104.8 16.545 104.975 17.425 ;
      RECT 104.8 16.915 107.425 17.085 ;
      RECT 103.475 16.545 104.975 16.715 ;
      RECT 104.315 15.695 104.645 16.715 ;
      RECT 103.475 15.695 103.805 16.715 ;
      RECT 102.455 22.775 102.785 23.295 ;
      RECT 102.665 22.025 102.835 22.86 ;
      RECT 102.61 22.735 102.835 22.86 ;
      RECT 102.62 22.025 102.835 22.155 ;
      RECT 102.445 21.18 102.775 22.105 ;
      RECT 101.615 22.775 101.945 23.3 ;
      RECT 101.745 22.275 101.945 23.3 ;
      RECT 101.745 22.275 102.495 22.605 ;
      RECT 101.745 21.135 101.935 23.3 ;
      RECT 101.04 21.695 101.935 22.07 ;
      RECT 101.595 21.135 101.935 22.07 ;
      RECT 100.085 23.065 100.87 23.235 ;
      RECT 100.7 21.265 100.87 23.235 ;
      RECT 100.7 22.275 101.575 22.605 ;
      RECT 99.985 21.265 100.87 21.435 ;
      RECT 97.575 11.815 97.745 12.465 ;
      RECT 98.415 11.815 98.585 12.46 ;
      RECT 97.575 11.815 98.995 11.985 ;
      RECT 98.82 11.105 98.995 11.985 ;
      RECT 98.82 11.475 101.445 11.645 ;
      RECT 97.495 11.105 98.995 11.275 ;
      RECT 98.335 10.255 98.665 11.275 ;
      RECT 97.495 10.255 97.825 11.275 ;
      RECT 100.605 19.655 100.935 20.58 ;
      RECT 100.825 18.9 100.995 19.735 ;
      RECT 100.78 19.605 100.995 19.735 ;
      RECT 100.77 18.9 100.995 19.025 ;
      RECT 100.615 18.465 100.945 18.985 ;
      RECT 99.755 19.69 100.095 20.625 ;
      RECT 99.905 18.46 100.095 20.625 ;
      RECT 99.2 19.69 100.095 20.065 ;
      RECT 99.905 19.155 100.655 19.485 ;
      RECT 99.905 18.46 100.105 19.485 ;
      RECT 99.775 18.46 100.105 18.985 ;
      RECT 100.065 22.565 100.53 22.895 ;
      RECT 100.21 21.605 100.53 22.895 ;
      RECT 99.51 23.065 99.915 23.235 ;
      RECT 99.51 21.135 99.68 23.235 ;
      RECT 98.85 22.535 99.68 22.835 ;
      RECT 98.85 22.505 99.05 22.835 ;
      RECT 99.51 21.135 99.76 21.465 ;
      RECT 98.145 20.325 99.03 20.495 ;
      RECT 98.86 18.525 99.03 20.495 ;
      RECT 98.86 19.155 99.735 19.485 ;
      RECT 98.245 18.525 99.03 18.695 ;
      RECT 97.965 23.065 98.64 23.235 ;
      RECT 98.47 22.115 98.64 23.235 ;
      RECT 99.17 22.025 99.34 22.355 ;
      RECT 98.47 22.115 99.34 22.285 ;
      RECT 98.83 22.025 99.34 22.285 ;
      RECT 98.83 21.24 99 22.285 ;
      RECT 97.895 21.24 99 21.41 ;
      RECT 98.37 18.865 98.69 20.155 ;
      RECT 98.225 18.865 98.69 19.195 ;
      RECT 97.775 22.645 98.3 22.865 ;
      RECT 98.13 21.58 98.3 22.865 ;
      RECT 98.13 21.58 98.66 21.945 ;
      RECT 97.845 25.095 98.175 26.02 ;
      RECT 98.065 24.34 98.235 25.175 ;
      RECT 98.02 25.045 98.235 25.175 ;
      RECT 98.01 24.34 98.235 24.465 ;
      RECT 97.855 23.905 98.185 24.425 ;
      RECT 97.975 17.255 98.145 17.905 ;
      RECT 95.715 17.655 97.25 17.905 ;
      RECT 97.08 17.255 97.25 17.905 ;
      RECT 95.715 17.255 95.885 17.905 ;
      RECT 97.08 17.255 98.145 17.425 ;
      RECT 95.085 17.255 95.885 17.425 ;
      RECT 95.085 16.535 95.255 17.425 ;
      RECT 95.085 16.535 98.145 16.705 ;
      RECT 97.975 15.695 98.145 16.705 ;
      RECT 97.67 20.295 97.92 20.625 ;
      RECT 97.67 18.525 97.84 20.625 ;
      RECT 97.01 18.925 97.21 19.255 ;
      RECT 97.01 18.925 97.84 19.225 ;
      RECT 97.67 18.525 98.075 18.695 ;
      RECT 96.995 25.13 97.335 26.065 ;
      RECT 97.145 23.9 97.335 26.065 ;
      RECT 96.44 25.13 97.335 25.505 ;
      RECT 97.145 24.595 97.895 24.925 ;
      RECT 97.145 23.9 97.345 24.925 ;
      RECT 97.015 23.9 97.345 24.425 ;
      RECT 97.475 15.695 97.805 16.365 ;
      RECT 96.635 15.695 96.965 15.905 ;
      RECT 96.635 15.695 97.805 15.865 ;
      RECT 97.435 23.065 97.77 23.235 ;
      RECT 97.435 22.795 97.605 23.235 ;
      RECT 97.38 21.56 97.55 22.925 ;
      RECT 97.435 21.135 97.685 21.69 ;
      RECT 96.055 20.35 97.16 20.52 ;
      RECT 96.99 19.475 97.16 20.52 ;
      RECT 96.99 19.475 97.5 19.735 ;
      RECT 97.33 19.405 97.5 19.735 ;
      RECT 96.63 19.475 97.5 19.645 ;
      RECT 96.63 18.525 96.8 19.645 ;
      RECT 96.125 18.525 96.8 18.695 ;
      RECT 95.67 16.125 97.305 16.365 ;
      RECT 97.075 16.035 97.305 16.365 ;
      RECT 95.67 15.695 95.92 16.365 ;
      RECT 97.04 30.835 97.295 31.505 ;
      RECT 97.125 29.295 97.295 31.505 ;
      RECT 97.11 29.295 97.295 29.705 ;
      RECT 97.085 29.295 97.295 29.635 ;
      RECT 97.04 29.295 97.295 29.625 ;
      RECT 96.62 16.885 96.9 17.485 ;
      RECT 96.62 16.885 97.095 17.085 ;
      RECT 95.385 25.765 96.27 25.935 ;
      RECT 96.1 23.965 96.27 25.935 ;
      RECT 96.1 24.595 96.975 24.925 ;
      RECT 95.485 23.965 96.27 24.135 ;
      RECT 93.895 30.495 94.065 31.505 ;
      RECT 93.895 30.495 96.955 30.665 ;
      RECT 96.785 29.775 96.955 30.665 ;
      RECT 96.155 29.775 96.955 29.945 ;
      RECT 93.895 29.775 94.96 29.945 ;
      RECT 94.79 29.295 94.96 29.945 ;
      RECT 96.155 29.295 96.325 29.945 ;
      RECT 93.895 29.295 94.065 29.945 ;
      RECT 94.79 29.295 96.325 29.545 ;
      RECT 96.29 19.815 96.82 20.18 ;
      RECT 96.29 18.895 96.46 20.18 ;
      RECT 95.935 18.895 96.46 19.115 ;
      RECT 96.19 30.145 96.565 30.315 ;
      RECT 96.19 30.115 96.555 30.315 ;
      RECT 95.735 22.795 95.905 23.255 ;
      RECT 95.735 22.795 96.4 22.965 ;
      RECT 96.17 21.635 96.4 22.965 ;
      RECT 95.735 21.635 96.4 21.805 ;
      RECT 95.735 21.135 95.905 21.805 ;
      RECT 96.12 14.515 96.375 15.185 ;
      RECT 96.205 12.975 96.375 15.185 ;
      RECT 96.19 12.975 96.375 13.385 ;
      RECT 96.16 12.975 96.375 13.315 ;
      RECT 96.12 12.975 96.375 13.305 ;
      RECT 96.12 30.835 96.37 31.505 ;
      RECT 94.735 30.835 94.965 31.165 ;
      RECT 94.735 30.835 96.37 31.075 ;
      RECT 96.065 16.885 96.35 17.485 ;
      RECT 96.02 16.885 96.35 17.085 ;
      RECT 92.975 14.175 93.145 15.185 ;
      RECT 92.975 14.175 96.035 14.345 ;
      RECT 95.865 13.455 96.035 14.345 ;
      RECT 95.235 13.455 96.035 13.625 ;
      RECT 92.975 13.455 94.04 13.625 ;
      RECT 93.87 12.975 94.04 13.625 ;
      RECT 95.235 12.975 95.405 13.625 ;
      RECT 92.975 12.975 93.145 13.625 ;
      RECT 93.87 12.975 95.405 13.225 ;
      RECT 95.69 30.115 96.02 30.315 ;
      RECT 95.69 29.715 95.975 30.315 ;
      RECT 95.595 20.07 95.845 20.625 ;
      RECT 95.54 18.835 95.71 20.2 ;
      RECT 95.595 18.525 95.765 18.965 ;
      RECT 95.595 18.525 95.93 18.695 ;
      RECT 95.61 24.305 95.93 25.595 ;
      RECT 95.465 24.305 95.93 24.635 ;
      RECT 95.485 16.885 95.85 17.085 ;
      RECT 95.475 16.885 95.85 17.055 ;
      RECT 95.27 13.825 95.645 13.995 ;
      RECT 95.27 13.795 95.635 13.995 ;
      RECT 91.595 11.815 91.765 12.465 ;
      RECT 92.435 11.815 92.605 12.46 ;
      RECT 91.595 11.815 93.015 11.985 ;
      RECT 92.84 11.105 93.015 11.985 ;
      RECT 92.84 11.475 95.465 11.645 ;
      RECT 91.515 11.105 93.015 11.275 ;
      RECT 92.355 10.255 92.685 11.275 ;
      RECT 91.515 10.255 91.845 11.275 ;
      RECT 95.2 14.515 95.45 15.185 ;
      RECT 93.815 14.515 94.045 14.845 ;
      RECT 93.815 14.515 95.45 14.755 ;
      RECT 94.945 30.115 95.42 30.315 ;
      RECT 95.14 29.715 95.42 30.315 ;
      RECT 94.235 31.335 95.405 31.505 ;
      RECT 95.075 31.295 95.405 31.505 ;
      RECT 94.235 30.835 94.565 31.505 ;
      RECT 94.91 25.735 95.16 26.065 ;
      RECT 94.91 23.965 95.08 26.065 ;
      RECT 94.25 24.365 94.45 24.695 ;
      RECT 94.25 24.365 95.08 24.665 ;
      RECT 94.91 23.965 95.315 24.135 ;
      RECT 94.77 13.795 95.1 13.995 ;
      RECT 94.77 13.395 95.055 13.995 ;
      RECT 94.745 17.575 95 17.905 ;
      RECT 94.745 17.565 94.955 17.905 ;
      RECT 94.745 17.495 94.93 17.905 ;
      RECT 94.745 15.695 94.915 17.905 ;
      RECT 94.745 15.695 95 16.365 ;
      RECT 93.295 25.79 94.4 25.96 ;
      RECT 94.23 24.915 94.4 25.96 ;
      RECT 94.23 24.915 94.74 25.175 ;
      RECT 94.57 24.845 94.74 25.175 ;
      RECT 93.87 24.915 94.74 25.085 ;
      RECT 93.87 23.965 94.04 25.085 ;
      RECT 93.365 23.965 94.04 24.135 ;
      RECT 93.895 19.955 94.065 20.625 ;
      RECT 93.895 19.955 94.56 20.125 ;
      RECT 94.33 18.795 94.56 20.125 ;
      RECT 93.895 18.795 94.56 18.965 ;
      RECT 93.895 18.505 94.065 18.965 ;
      RECT 94.025 13.795 94.5 13.995 ;
      RECT 94.22 13.395 94.5 13.995 ;
      RECT 93.315 15.015 94.485 15.185 ;
      RECT 94.155 14.975 94.485 15.185 ;
      RECT 93.315 14.515 93.645 15.185 ;
      RECT 93.53 25.255 94.06 25.62 ;
      RECT 93.53 24.335 93.7 25.62 ;
      RECT 93.175 24.335 93.7 24.555 ;
      RECT 92.835 25.51 93.085 26.065 ;
      RECT 92.78 24.275 92.95 25.64 ;
      RECT 92.835 23.965 93.005 24.405 ;
      RECT 92.835 23.965 93.17 24.135 ;
      RECT 91.135 25.395 91.305 26.065 ;
      RECT 91.135 25.395 91.8 25.565 ;
      RECT 91.57 24.235 91.8 25.565 ;
      RECT 91.135 24.235 91.8 24.405 ;
      RECT 91.135 23.945 91.305 24.405 ;
      RECT 87.735 22.775 88.065 23.295 ;
      RECT 87.945 22.025 88.115 22.86 ;
      RECT 87.89 22.735 88.115 22.86 ;
      RECT 87.9 22.025 88.115 22.155 ;
      RECT 87.725 21.18 88.055 22.105 ;
      RECT 86.895 22.775 87.225 23.3 ;
      RECT 87.025 22.275 87.225 23.3 ;
      RECT 87.025 22.275 87.775 22.605 ;
      RECT 87.025 21.135 87.215 23.3 ;
      RECT 86.32 21.695 87.215 22.07 ;
      RECT 86.875 21.135 87.215 22.07 ;
      RECT 85.365 23.065 86.15 23.235 ;
      RECT 85.98 21.265 86.15 23.235 ;
      RECT 85.98 22.275 86.855 22.605 ;
      RECT 85.265 21.265 86.15 21.435 ;
      RECT 82.855 11.815 83.025 12.465 ;
      RECT 83.695 11.815 83.865 12.46 ;
      RECT 82.855 11.815 84.275 11.985 ;
      RECT 84.1 11.105 84.275 11.985 ;
      RECT 84.1 11.475 86.725 11.645 ;
      RECT 82.775 11.105 84.275 11.275 ;
      RECT 83.615 10.255 83.945 11.275 ;
      RECT 82.775 10.255 83.105 11.275 ;
      RECT 86 19.955 86.255 20.625 ;
      RECT 86.085 18.415 86.255 20.625 ;
      RECT 86.07 18.415 86.255 18.825 ;
      RECT 86 18.415 86.255 18.745 ;
      RECT 82.855 19.615 83.025 20.625 ;
      RECT 82.855 19.615 85.915 19.785 ;
      RECT 85.745 18.895 85.915 19.785 ;
      RECT 85.115 18.895 85.915 19.065 ;
      RECT 82.855 18.895 83.92 19.065 ;
      RECT 83.75 18.415 83.92 19.065 ;
      RECT 85.115 18.415 85.285 19.065 ;
      RECT 82.855 18.415 83.025 19.065 ;
      RECT 83.75 18.415 85.285 18.665 ;
      RECT 85.345 22.565 85.81 22.895 ;
      RECT 85.49 21.605 85.81 22.895 ;
      RECT 85.15 19.265 85.525 19.435 ;
      RECT 85.15 19.235 85.515 19.435 ;
      RECT 85.08 19.955 85.33 20.625 ;
      RECT 83.695 19.955 83.925 20.285 ;
      RECT 83.695 19.955 85.33 20.195 ;
      RECT 84.79 23.065 85.195 23.235 ;
      RECT 84.79 21.135 84.96 23.235 ;
      RECT 84.13 22.535 84.96 22.835 ;
      RECT 84.13 22.505 84.33 22.835 ;
      RECT 84.79 21.135 85.04 21.465 ;
      RECT 84.65 19.235 84.98 19.435 ;
      RECT 84.65 18.835 84.935 19.435 ;
      RECT 84.635 17.255 84.805 17.905 ;
      RECT 82.375 17.655 83.91 17.905 ;
      RECT 83.74 17.255 83.91 17.905 ;
      RECT 82.375 17.255 82.545 17.905 ;
      RECT 83.74 17.255 84.805 17.425 ;
      RECT 81.745 17.255 82.545 17.425 ;
      RECT 81.745 16.535 81.915 17.425 ;
      RECT 81.745 16.535 84.805 16.705 ;
      RECT 84.635 15.695 84.805 16.705 ;
      RECT 83.245 23.065 83.92 23.235 ;
      RECT 83.75 22.115 83.92 23.235 ;
      RECT 84.45 22.025 84.62 22.355 ;
      RECT 83.75 22.115 84.62 22.285 ;
      RECT 84.11 22.025 84.62 22.285 ;
      RECT 84.11 21.24 84.28 22.285 ;
      RECT 83.175 21.24 84.28 21.41 ;
      RECT 84.135 15.695 84.465 16.365 ;
      RECT 83.295 15.695 83.625 15.905 ;
      RECT 83.295 15.695 84.465 15.865 ;
      RECT 84.045 25.095 84.375 26.02 ;
      RECT 84.265 24.34 84.435 25.175 ;
      RECT 84.22 25.045 84.435 25.175 ;
      RECT 84.21 24.34 84.435 24.465 ;
      RECT 84.055 23.905 84.385 24.425 ;
      RECT 83.905 19.235 84.38 19.435 ;
      RECT 84.1 18.835 84.38 19.435 ;
      RECT 83.195 20.455 84.365 20.625 ;
      RECT 84.035 20.415 84.365 20.625 ;
      RECT 83.195 19.955 83.525 20.625 ;
      RECT 83.195 25.13 83.535 26.065 ;
      RECT 83.345 23.9 83.535 26.065 ;
      RECT 82.64 25.13 83.535 25.505 ;
      RECT 83.345 24.595 84.095 24.925 ;
      RECT 83.345 23.9 83.545 24.925 ;
      RECT 83.215 23.9 83.545 24.425 ;
      RECT 82.33 16.125 83.965 16.365 ;
      RECT 83.735 16.035 83.965 16.365 ;
      RECT 82.33 15.695 82.58 16.365 ;
      RECT 83.7 30.835 83.955 31.505 ;
      RECT 83.785 29.295 83.955 31.505 ;
      RECT 83.77 29.295 83.955 29.705 ;
      RECT 83.745 29.295 83.955 29.635 ;
      RECT 83.7 29.295 83.955 29.625 ;
      RECT 83.055 22.645 83.58 22.865 ;
      RECT 83.41 21.58 83.58 22.865 ;
      RECT 83.41 21.58 83.94 21.945 ;
      RECT 83.28 16.885 83.56 17.485 ;
      RECT 83.28 16.885 83.755 17.085 ;
      RECT 80.555 30.495 80.725 31.505 ;
      RECT 80.555 30.495 83.615 30.665 ;
      RECT 83.445 29.775 83.615 30.665 ;
      RECT 82.815 29.775 83.615 29.945 ;
      RECT 80.555 29.775 81.62 29.945 ;
      RECT 81.45 29.295 81.62 29.945 ;
      RECT 82.815 29.295 82.985 29.945 ;
      RECT 80.555 29.295 80.725 29.945 ;
      RECT 81.45 29.295 82.985 29.545 ;
      RECT 82.85 30.145 83.225 30.315 ;
      RECT 82.85 30.115 83.215 30.315 ;
      RECT 81.585 25.765 82.47 25.935 ;
      RECT 82.3 23.965 82.47 25.935 ;
      RECT 82.3 24.595 83.175 24.925 ;
      RECT 81.685 23.965 82.47 24.135 ;
      RECT 82.715 23.065 83.05 23.235 ;
      RECT 82.715 22.795 82.885 23.235 ;
      RECT 82.66 21.56 82.83 22.925 ;
      RECT 82.715 21.135 82.965 21.69 ;
      RECT 82.78 30.835 83.03 31.505 ;
      RECT 81.395 30.835 81.625 31.165 ;
      RECT 81.395 30.835 83.03 31.075 ;
      RECT 82.725 16.885 83.01 17.485 ;
      RECT 82.68 16.885 83.01 17.085 ;
      RECT 82.35 30.115 82.68 30.315 ;
      RECT 82.35 29.715 82.635 30.315 ;
      RECT 82.205 19.655 82.535 20.58 ;
      RECT 82.425 18.9 82.595 19.735 ;
      RECT 82.38 19.605 82.595 19.735 ;
      RECT 82.37 18.9 82.595 19.025 ;
      RECT 82.215 18.465 82.545 18.985 ;
      RECT 82.145 16.885 82.51 17.085 ;
      RECT 82.135 16.885 82.51 17.055 ;
      RECT 81.355 19.69 81.695 20.625 ;
      RECT 81.505 18.46 81.695 20.625 ;
      RECT 80.8 19.69 81.695 20.065 ;
      RECT 81.505 19.155 82.255 19.485 ;
      RECT 81.505 18.46 81.705 19.485 ;
      RECT 81.375 18.46 81.705 18.985 ;
      RECT 81.81 24.305 82.13 25.595 ;
      RECT 81.665 24.305 82.13 24.635 ;
      RECT 81.605 30.115 82.08 30.315 ;
      RECT 81.8 29.715 82.08 30.315 ;
      RECT 80.895 31.335 82.065 31.505 ;
      RECT 81.735 31.295 82.065 31.505 ;
      RECT 80.895 30.835 81.225 31.505 ;
      RECT 81.015 22.795 81.185 23.255 ;
      RECT 81.015 22.795 81.68 22.965 ;
      RECT 81.45 21.635 81.68 22.965 ;
      RECT 81.015 21.635 81.68 21.805 ;
      RECT 81.015 21.135 81.185 21.805 ;
      RECT 81.405 17.575 81.66 17.905 ;
      RECT 81.405 17.565 81.615 17.905 ;
      RECT 81.405 17.495 81.59 17.905 ;
      RECT 81.405 15.695 81.575 17.905 ;
      RECT 81.405 15.695 81.66 16.365 ;
      RECT 81.11 25.735 81.36 26.065 ;
      RECT 81.11 23.965 81.28 26.065 ;
      RECT 80.45 24.365 80.65 24.695 ;
      RECT 80.45 24.365 81.28 24.665 ;
      RECT 81.11 23.965 81.515 24.135 ;
      RECT 79.745 20.325 80.63 20.495 ;
      RECT 80.46 18.525 80.63 20.495 ;
      RECT 80.46 19.155 81.335 19.485 ;
      RECT 79.845 18.525 80.63 18.695 ;
      RECT 79.495 25.79 80.6 25.96 ;
      RECT 80.43 24.915 80.6 25.96 ;
      RECT 80.43 24.915 80.94 25.175 ;
      RECT 80.77 24.845 80.94 25.175 ;
      RECT 80.07 24.915 80.94 25.085 ;
      RECT 80.07 23.965 80.24 25.085 ;
      RECT 79.565 23.965 80.24 24.135 ;
      RECT 80.495 22.84 80.755 23.345 ;
      RECT 80.585 21.135 80.755 23.345 ;
      RECT 80.485 21.135 80.755 22.04 ;
      RECT 79.635 22.795 79.805 23.345 ;
      RECT 79.635 22.795 80.3 22.965 ;
      RECT 80.13 21.895 80.3 22.965 ;
      RECT 80.13 22.21 80.415 22.54 ;
      RECT 79.635 21.895 80.3 22.065 ;
      RECT 79.635 21.135 79.805 22.065 ;
      RECT 79.97 18.865 80.29 20.155 ;
      RECT 79.825 18.865 80.29 19.195 ;
      RECT 79.73 25.255 80.26 25.62 ;
      RECT 79.73 24.335 79.9 25.62 ;
      RECT 79.375 24.335 79.9 24.555 ;
      RECT 79.27 20.295 79.52 20.625 ;
      RECT 79.27 18.525 79.44 20.625 ;
      RECT 78.61 18.925 78.81 19.255 ;
      RECT 78.61 18.925 79.44 19.225 ;
      RECT 79.27 18.525 79.675 18.695 ;
      RECT 79.035 25.51 79.285 26.065 ;
      RECT 78.98 24.275 79.15 25.64 ;
      RECT 79.035 23.965 79.205 24.405 ;
      RECT 79.035 23.965 79.37 24.135 ;
      RECT 77.655 20.35 78.76 20.52 ;
      RECT 78.59 19.475 78.76 20.52 ;
      RECT 78.59 19.475 79.1 19.735 ;
      RECT 78.93 19.405 79.1 19.735 ;
      RECT 78.23 19.475 79.1 19.645 ;
      RECT 78.23 18.525 78.4 19.645 ;
      RECT 77.725 18.525 78.4 18.695 ;
      RECT 77.89 19.815 78.42 20.18 ;
      RECT 77.89 18.895 78.06 20.18 ;
      RECT 77.535 18.895 78.06 19.115 ;
      RECT 77.335 25.395 77.505 26.065 ;
      RECT 77.335 25.395 78 25.565 ;
      RECT 77.77 24.235 78 25.565 ;
      RECT 77.335 24.235 78 24.405 ;
      RECT 77.335 23.945 77.505 24.405 ;
      RECT 74.115 11.815 74.285 12.465 ;
      RECT 74.955 11.815 75.125 12.46 ;
      RECT 74.115 11.815 75.535 11.985 ;
      RECT 75.36 11.105 75.535 11.985 ;
      RECT 75.36 11.475 77.985 11.645 ;
      RECT 74.035 11.105 75.535 11.275 ;
      RECT 74.875 10.255 75.205 11.275 ;
      RECT 74.035 10.255 74.365 11.275 ;
      RECT 74.115 17.255 74.285 17.905 ;
      RECT 74.955 17.255 75.125 17.9 ;
      RECT 74.115 17.255 75.535 17.425 ;
      RECT 75.36 16.545 75.535 17.425 ;
      RECT 75.36 16.915 77.985 17.085 ;
      RECT 74.035 16.545 75.535 16.715 ;
      RECT 74.875 15.695 75.205 16.715 ;
      RECT 74.035 15.695 74.365 16.715 ;
      RECT 77.195 20.07 77.445 20.625 ;
      RECT 77.14 18.835 77.31 20.2 ;
      RECT 77.195 18.525 77.365 18.965 ;
      RECT 77.195 18.525 77.53 18.695 ;
      RECT 77.26 30.835 77.515 31.505 ;
      RECT 77.345 29.295 77.515 31.505 ;
      RECT 77.33 29.295 77.515 29.705 ;
      RECT 77.305 29.295 77.515 29.635 ;
      RECT 77.26 29.295 77.515 29.625 ;
      RECT 74.115 30.495 74.285 31.505 ;
      RECT 74.115 30.495 77.175 30.665 ;
      RECT 77.005 29.775 77.175 30.665 ;
      RECT 76.375 29.775 77.175 29.945 ;
      RECT 74.115 29.775 75.18 29.945 ;
      RECT 75.01 29.295 75.18 29.945 ;
      RECT 76.375 29.295 76.545 29.945 ;
      RECT 74.115 29.295 74.285 29.945 ;
      RECT 75.01 29.295 76.545 29.545 ;
      RECT 76.41 30.145 76.785 30.315 ;
      RECT 76.41 30.115 76.775 30.315 ;
      RECT 76.34 30.835 76.59 31.505 ;
      RECT 74.955 30.835 75.185 31.165 ;
      RECT 74.955 30.835 76.59 31.075 ;
      RECT 75.91 30.115 76.24 30.315 ;
      RECT 75.91 29.715 76.195 30.315 ;
      RECT 75.495 19.955 75.665 20.625 ;
      RECT 75.495 19.955 76.16 20.125 ;
      RECT 75.93 18.795 76.16 20.125 ;
      RECT 75.495 18.795 76.16 18.965 ;
      RECT 75.495 18.505 75.665 18.965 ;
      RECT 75.165 30.115 75.64 30.315 ;
      RECT 75.36 29.715 75.64 30.315 ;
      RECT 74.455 31.335 75.625 31.505 ;
      RECT 75.295 31.295 75.625 31.505 ;
      RECT 74.455 30.835 74.785 31.505 ;
      RECT 73.015 22.775 73.345 23.295 ;
      RECT 73.225 22.025 73.395 22.86 ;
      RECT 73.17 22.735 73.395 22.86 ;
      RECT 73.18 22.025 73.395 22.155 ;
      RECT 73.005 21.18 73.335 22.105 ;
      RECT 72.175 22.775 72.505 23.3 ;
      RECT 72.305 22.275 72.505 23.3 ;
      RECT 72.305 22.275 73.055 22.605 ;
      RECT 72.305 21.135 72.495 23.3 ;
      RECT 71.6 21.695 72.495 22.07 ;
      RECT 72.155 21.135 72.495 22.07 ;
      RECT 70.645 23.065 71.43 23.235 ;
      RECT 71.26 21.265 71.43 23.235 ;
      RECT 71.26 22.275 72.135 22.605 ;
      RECT 70.545 21.265 71.43 21.435 ;
      RECT 71.755 17.255 71.925 17.905 ;
      RECT 69.495 17.655 71.03 17.905 ;
      RECT 70.86 17.255 71.03 17.905 ;
      RECT 69.495 17.255 69.665 17.905 ;
      RECT 70.86 17.255 71.925 17.425 ;
      RECT 68.865 17.255 69.665 17.425 ;
      RECT 68.865 16.535 69.035 17.425 ;
      RECT 68.865 16.535 71.925 16.705 ;
      RECT 71.755 15.695 71.925 16.705 ;
      RECT 71.755 19.615 71.925 20.625 ;
      RECT 68.865 19.615 71.925 19.785 ;
      RECT 68.865 18.895 69.035 19.785 ;
      RECT 70.86 18.895 71.925 19.065 ;
      RECT 71.755 18.415 71.925 19.065 ;
      RECT 68.865 18.895 69.665 19.065 ;
      RECT 69.495 18.415 69.665 19.065 ;
      RECT 70.86 18.415 71.03 19.065 ;
      RECT 69.495 18.415 71.03 18.665 ;
      RECT 71.755 28.135 71.925 28.785 ;
      RECT 69.495 28.535 71.03 28.785 ;
      RECT 70.86 28.135 71.03 28.785 ;
      RECT 69.495 28.135 69.665 28.785 ;
      RECT 70.86 28.135 71.925 28.305 ;
      RECT 68.865 28.135 69.665 28.305 ;
      RECT 68.865 27.415 69.035 28.305 ;
      RECT 68.865 27.415 71.925 27.585 ;
      RECT 71.755 26.575 71.925 27.585 ;
      RECT 71.255 15.695 71.585 16.365 ;
      RECT 70.415 15.695 70.745 15.905 ;
      RECT 70.415 15.695 71.585 15.865 ;
      RECT 70.415 20.455 71.585 20.625 ;
      RECT 71.255 19.955 71.585 20.625 ;
      RECT 70.415 20.415 70.745 20.625 ;
      RECT 71.255 26.575 71.585 27.245 ;
      RECT 70.415 26.575 70.745 26.785 ;
      RECT 70.415 26.575 71.585 26.745 ;
      RECT 70.625 22.565 71.09 22.895 ;
      RECT 70.77 21.605 71.09 22.895 ;
      RECT 69.45 16.125 71.085 16.365 ;
      RECT 70.855 16.035 71.085 16.365 ;
      RECT 69.45 15.695 69.7 16.365 ;
      RECT 69.45 19.955 69.7 20.625 ;
      RECT 70.855 19.955 71.085 20.285 ;
      RECT 69.45 19.955 71.085 20.195 ;
      RECT 69.45 27.005 71.085 27.245 ;
      RECT 70.855 26.915 71.085 27.245 ;
      RECT 69.45 26.575 69.7 27.245 ;
      RECT 70.4 16.885 70.68 17.485 ;
      RECT 70.4 16.885 70.875 17.085 ;
      RECT 70.4 19.235 70.875 19.435 ;
      RECT 70.4 18.835 70.68 19.435 ;
      RECT 70.4 27.765 70.68 28.365 ;
      RECT 70.4 27.765 70.875 27.965 ;
      RECT 70.07 23.065 70.475 23.235 ;
      RECT 70.07 21.135 70.24 23.235 ;
      RECT 69.41 22.535 70.24 22.835 ;
      RECT 69.41 22.505 69.61 22.835 ;
      RECT 70.07 21.135 70.32 21.465 ;
      RECT 69.845 16.885 70.13 17.485 ;
      RECT 69.8 16.885 70.13 17.085 ;
      RECT 69.8 19.235 70.13 19.435 ;
      RECT 69.845 18.835 70.13 19.435 ;
      RECT 69.845 27.765 70.13 28.365 ;
      RECT 69.8 27.765 70.13 27.965 ;
      RECT 68.525 23.065 69.2 23.235 ;
      RECT 69.03 22.115 69.2 23.235 ;
      RECT 69.73 22.025 69.9 22.355 ;
      RECT 69.03 22.115 69.9 22.285 ;
      RECT 69.39 22.025 69.9 22.285 ;
      RECT 69.39 21.24 69.56 22.285 ;
      RECT 68.455 21.24 69.56 21.41 ;
      RECT 66.595 14.165 66.925 15.185 ;
      RECT 65.755 14.165 66.085 15.185 ;
      RECT 65.755 14.165 67.255 14.335 ;
      RECT 67.08 13.455 67.255 14.335 ;
      RECT 67.08 13.795 69.705 13.965 ;
      RECT 65.835 13.455 67.255 13.625 ;
      RECT 66.675 12.98 66.845 13.625 ;
      RECT 65.835 12.975 66.005 13.625 ;
      RECT 66.595 25.045 66.925 26.065 ;
      RECT 65.755 25.045 66.085 26.065 ;
      RECT 65.755 25.045 67.255 25.215 ;
      RECT 67.08 24.335 67.255 25.215 ;
      RECT 67.08 24.675 69.705 24.845 ;
      RECT 65.835 24.335 67.255 24.505 ;
      RECT 66.675 23.86 66.845 24.505 ;
      RECT 65.835 23.855 66.005 24.505 ;
      RECT 69.265 16.885 69.63 17.085 ;
      RECT 69.255 16.885 69.63 17.055 ;
      RECT 69.255 19.265 69.63 19.435 ;
      RECT 69.265 19.235 69.63 19.435 ;
      RECT 69.265 27.765 69.63 27.965 ;
      RECT 69.255 27.765 69.63 27.935 ;
      RECT 68.335 22.645 68.86 22.865 ;
      RECT 68.69 21.58 68.86 22.865 ;
      RECT 68.69 21.58 69.22 21.945 ;
      RECT 68.525 17.575 68.78 17.905 ;
      RECT 68.525 17.565 68.735 17.905 ;
      RECT 68.525 17.495 68.71 17.905 ;
      RECT 68.525 15.695 68.695 17.905 ;
      RECT 68.525 15.695 68.78 16.365 ;
      RECT 68.525 19.955 68.78 20.625 ;
      RECT 68.525 18.415 68.695 20.625 ;
      RECT 68.525 18.415 68.71 18.825 ;
      RECT 68.525 18.415 68.78 18.745 ;
      RECT 68.525 28.455 68.78 28.785 ;
      RECT 68.525 28.445 68.735 28.785 ;
      RECT 68.525 28.375 68.71 28.785 ;
      RECT 68.525 26.575 68.695 28.785 ;
      RECT 68.525 26.575 68.78 27.245 ;
      RECT 67.995 23.065 68.33 23.235 ;
      RECT 67.995 22.795 68.165 23.235 ;
      RECT 67.94 21.56 68.11 22.925 ;
      RECT 67.995 21.135 68.245 21.69 ;
      RECT 66.295 22.795 66.465 23.255 ;
      RECT 66.295 22.795 66.96 22.965 ;
      RECT 66.73 21.635 66.96 22.965 ;
      RECT 66.295 21.635 66.96 21.805 ;
      RECT 66.295 21.135 66.465 21.805 ;
      RECT 66.115 17.335 66.445 17.855 ;
      RECT 66.325 16.585 66.495 17.42 ;
      RECT 66.27 17.295 66.495 17.42 ;
      RECT 66.28 16.585 66.495 16.715 ;
      RECT 66.105 15.74 66.435 16.665 ;
      RECT 66.105 19.655 66.435 20.58 ;
      RECT 66.325 18.9 66.495 19.735 ;
      RECT 66.28 19.605 66.495 19.735 ;
      RECT 66.27 18.9 66.495 19.025 ;
      RECT 66.115 18.465 66.445 18.985 ;
      RECT 66.115 28.215 66.445 28.735 ;
      RECT 66.325 27.465 66.495 28.3 ;
      RECT 66.27 28.175 66.495 28.3 ;
      RECT 66.28 27.465 66.495 27.595 ;
      RECT 66.105 26.62 66.435 27.545 ;
      RECT 66.105 30.535 66.435 31.46 ;
      RECT 66.325 29.78 66.495 30.615 ;
      RECT 66.28 30.485 66.495 30.615 ;
      RECT 66.27 29.78 66.495 29.905 ;
      RECT 66.115 29.345 66.445 29.865 ;
      RECT 62.615 11.815 62.785 12.465 ;
      RECT 63.455 11.815 63.625 12.46 ;
      RECT 62.615 11.815 64.035 11.985 ;
      RECT 63.86 11.105 64.035 11.985 ;
      RECT 63.86 11.475 66.485 11.645 ;
      RECT 62.535 11.105 64.035 11.275 ;
      RECT 63.375 10.255 63.705 11.275 ;
      RECT 62.535 10.255 62.865 11.275 ;
      RECT 65.275 17.335 65.605 17.86 ;
      RECT 65.405 16.835 65.605 17.86 ;
      RECT 65.405 16.835 66.155 17.165 ;
      RECT 65.405 15.695 65.595 17.86 ;
      RECT 64.7 16.255 65.595 16.63 ;
      RECT 65.255 15.695 65.595 16.63 ;
      RECT 65.255 19.69 65.595 20.625 ;
      RECT 65.405 18.46 65.595 20.625 ;
      RECT 64.7 19.69 65.595 20.065 ;
      RECT 65.405 19.155 66.155 19.485 ;
      RECT 65.405 18.46 65.605 19.485 ;
      RECT 65.275 18.46 65.605 18.985 ;
      RECT 65.275 28.215 65.605 28.74 ;
      RECT 65.405 27.715 65.605 28.74 ;
      RECT 65.405 27.715 66.155 28.045 ;
      RECT 65.405 26.575 65.595 28.74 ;
      RECT 64.7 27.135 65.595 27.51 ;
      RECT 65.255 26.575 65.595 27.51 ;
      RECT 65.255 30.57 65.595 31.505 ;
      RECT 65.405 29.34 65.595 31.505 ;
      RECT 64.7 30.57 65.595 30.945 ;
      RECT 65.405 30.035 66.155 30.365 ;
      RECT 65.405 29.34 65.605 30.365 ;
      RECT 65.275 29.34 65.605 29.865 ;
      RECT 63.745 17.625 64.53 17.795 ;
      RECT 64.36 15.825 64.53 17.795 ;
      RECT 64.36 16.835 65.235 17.165 ;
      RECT 63.645 15.825 64.53 15.995 ;
      RECT 63.645 20.325 64.53 20.495 ;
      RECT 64.36 18.525 64.53 20.495 ;
      RECT 64.36 19.155 65.235 19.485 ;
      RECT 63.745 18.525 64.53 18.695 ;
      RECT 63.745 28.505 64.53 28.675 ;
      RECT 64.36 26.705 64.53 28.675 ;
      RECT 64.36 27.715 65.235 28.045 ;
      RECT 63.645 26.705 64.53 26.875 ;
      RECT 63.645 31.205 64.53 31.375 ;
      RECT 64.36 29.405 64.53 31.375 ;
      RECT 64.36 30.035 65.235 30.365 ;
      RECT 63.745 29.405 64.53 29.575 ;
      RECT 63.725 17.125 64.19 17.455 ;
      RECT 63.87 16.165 64.19 17.455 ;
      RECT 63.87 18.865 64.19 20.155 ;
      RECT 63.725 18.865 64.19 19.195 ;
      RECT 63.725 28.005 64.19 28.335 ;
      RECT 63.87 27.045 64.19 28.335 ;
      RECT 63.87 29.745 64.19 31.035 ;
      RECT 63.725 29.745 64.19 30.075 ;
      RECT 63.935 14.175 64.105 15.185 ;
      RECT 61.045 14.175 64.105 14.345 ;
      RECT 61.045 13.455 61.215 14.345 ;
      RECT 63.04 13.455 64.105 13.625 ;
      RECT 63.935 12.975 64.105 13.625 ;
      RECT 61.045 13.455 61.845 13.625 ;
      RECT 61.675 12.975 61.845 13.625 ;
      RECT 63.04 12.975 63.21 13.625 ;
      RECT 61.675 12.975 63.21 13.225 ;
      RECT 62.595 15.015 63.765 15.185 ;
      RECT 63.435 14.515 63.765 15.185 ;
      RECT 62.595 14.975 62.925 15.185 ;
      RECT 63.17 17.625 63.575 17.795 ;
      RECT 63.17 15.695 63.34 17.795 ;
      RECT 62.51 17.095 63.34 17.395 ;
      RECT 62.51 17.065 62.71 17.395 ;
      RECT 63.17 15.695 63.42 16.025 ;
      RECT 63.17 20.295 63.42 20.625 ;
      RECT 63.17 18.525 63.34 20.625 ;
      RECT 62.51 18.925 62.71 19.255 ;
      RECT 62.51 18.925 63.34 19.225 ;
      RECT 63.17 18.525 63.575 18.695 ;
      RECT 63.17 28.505 63.575 28.675 ;
      RECT 63.17 26.575 63.34 28.675 ;
      RECT 62.51 27.975 63.34 28.275 ;
      RECT 62.51 27.945 62.71 28.275 ;
      RECT 63.17 26.575 63.42 26.905 ;
      RECT 63.17 31.175 63.42 31.505 ;
      RECT 63.17 29.405 63.34 31.505 ;
      RECT 62.51 29.805 62.71 30.135 ;
      RECT 62.51 29.805 63.34 30.105 ;
      RECT 63.17 29.405 63.575 29.575 ;
      RECT 61.63 14.515 61.88 15.185 ;
      RECT 63.035 14.515 63.265 14.845 ;
      RECT 61.63 14.515 63.265 14.755 ;
      RECT 62.58 13.795 63.055 13.995 ;
      RECT 62.58 13.395 62.86 13.995 ;
      RECT 61.625 17.625 62.3 17.795 ;
      RECT 62.13 16.675 62.3 17.795 ;
      RECT 62.83 16.585 63 16.915 ;
      RECT 62.13 16.675 63 16.845 ;
      RECT 62.49 16.585 63 16.845 ;
      RECT 62.49 15.8 62.66 16.845 ;
      RECT 61.555 15.8 62.66 15.97 ;
      RECT 61.555 20.35 62.66 20.52 ;
      RECT 62.49 19.475 62.66 20.52 ;
      RECT 62.49 19.475 63 19.735 ;
      RECT 62.83 19.405 63 19.735 ;
      RECT 62.13 19.475 63 19.645 ;
      RECT 62.13 18.525 62.3 19.645 ;
      RECT 61.625 18.525 62.3 18.695 ;
      RECT 61.625 28.505 62.3 28.675 ;
      RECT 62.13 27.555 62.3 28.675 ;
      RECT 62.83 27.465 63 27.795 ;
      RECT 62.13 27.555 63 27.725 ;
      RECT 62.49 27.465 63 27.725 ;
      RECT 62.49 26.68 62.66 27.725 ;
      RECT 61.555 26.68 62.66 26.85 ;
      RECT 61.555 31.23 62.66 31.4 ;
      RECT 62.49 30.355 62.66 31.4 ;
      RECT 62.49 30.355 63 30.615 ;
      RECT 62.83 30.285 63 30.615 ;
      RECT 62.13 30.355 63 30.525 ;
      RECT 62.13 29.405 62.3 30.525 ;
      RECT 61.625 29.405 62.3 29.575 ;
      RECT 61.435 17.205 61.96 17.425 ;
      RECT 61.79 16.14 61.96 17.425 ;
      RECT 61.79 16.14 62.32 16.505 ;
      RECT 61.79 19.815 62.32 20.18 ;
      RECT 61.79 18.895 61.96 20.18 ;
      RECT 61.435 18.895 61.96 19.115 ;
      RECT 61.435 28.085 61.96 28.305 ;
      RECT 61.79 27.02 61.96 28.305 ;
      RECT 61.79 27.02 62.32 27.385 ;
      RECT 61.79 30.695 62.32 31.06 ;
      RECT 61.79 29.775 61.96 31.06 ;
      RECT 61.435 29.775 61.96 29.995 ;
      RECT 61.98 13.795 62.31 13.995 ;
      RECT 62.025 13.395 62.31 13.995 ;
      RECT 61.435 13.825 61.81 13.995 ;
      RECT 61.445 13.795 61.81 13.995 ;
      RECT 61.095 17.625 61.43 17.795 ;
      RECT 61.095 17.355 61.265 17.795 ;
      RECT 61.04 16.12 61.21 17.485 ;
      RECT 61.095 15.695 61.345 16.25 ;
      RECT 61.095 20.07 61.345 20.625 ;
      RECT 61.04 18.835 61.21 20.2 ;
      RECT 61.095 18.525 61.265 18.965 ;
      RECT 61.095 18.525 61.43 18.695 ;
      RECT 61.095 28.505 61.43 28.675 ;
      RECT 61.095 28.235 61.265 28.675 ;
      RECT 61.04 27 61.21 28.365 ;
      RECT 61.095 26.575 61.345 27.13 ;
      RECT 61.095 30.95 61.345 31.505 ;
      RECT 61.04 29.715 61.21 31.08 ;
      RECT 61.095 29.405 61.265 29.845 ;
      RECT 61.095 29.405 61.43 29.575 ;
      RECT 61.175 22.795 61.345 23.345 ;
      RECT 60.68 22.795 61.345 22.965 ;
      RECT 60.68 21.895 60.85 22.965 ;
      RECT 60.565 22.21 60.85 22.54 ;
      RECT 60.68 21.895 61.345 22.065 ;
      RECT 61.175 21.135 61.345 22.065 ;
      RECT 60.705 14.515 60.96 15.185 ;
      RECT 60.705 12.975 60.875 15.185 ;
      RECT 60.705 12.975 60.89 13.385 ;
      RECT 60.705 12.975 60.96 13.305 ;
      RECT 60.225 22.84 60.485 23.345 ;
      RECT 60.225 21.135 60.395 23.345 ;
      RECT 60.225 21.135 60.495 22.04 ;
      RECT 59.395 17.355 59.565 17.815 ;
      RECT 59.395 17.355 60.06 17.525 ;
      RECT 59.83 16.195 60.06 17.525 ;
      RECT 59.395 16.195 60.06 16.365 ;
      RECT 59.395 15.695 59.565 16.365 ;
      RECT 59.395 19.955 59.565 20.625 ;
      RECT 59.395 19.955 60.06 20.125 ;
      RECT 59.83 18.795 60.06 20.125 ;
      RECT 59.395 18.795 60.06 18.965 ;
      RECT 59.395 18.505 59.565 18.965 ;
      RECT 59.395 28.235 59.565 28.695 ;
      RECT 59.395 28.235 60.06 28.405 ;
      RECT 59.83 27.075 60.06 28.405 ;
      RECT 59.395 27.075 60.06 27.245 ;
      RECT 59.395 26.575 59.565 27.245 ;
      RECT 59.395 30.835 59.565 31.505 ;
      RECT 59.395 30.835 60.06 31.005 ;
      RECT 59.83 29.675 60.06 31.005 ;
      RECT 59.395 29.675 60.06 29.845 ;
      RECT 59.395 29.385 59.565 29.845 ;
      RECT 58.295 22.775 58.625 23.295 ;
      RECT 58.505 22.025 58.675 22.86 ;
      RECT 58.45 22.735 58.675 22.86 ;
      RECT 58.46 22.025 58.675 22.155 ;
      RECT 58.285 21.18 58.615 22.105 ;
      RECT 57.455 22.775 57.785 23.3 ;
      RECT 57.585 22.275 57.785 23.3 ;
      RECT 57.585 22.275 58.335 22.605 ;
      RECT 57.585 21.135 57.775 23.3 ;
      RECT 56.88 21.695 57.775 22.07 ;
      RECT 57.435 21.135 57.775 22.07 ;
      RECT 55.925 23.065 56.71 23.235 ;
      RECT 56.54 21.265 56.71 23.235 ;
      RECT 56.54 22.275 57.415 22.605 ;
      RECT 55.825 21.265 56.71 21.435 ;
      RECT 56.915 17.335 57.245 17.855 ;
      RECT 57.125 16.585 57.295 17.42 ;
      RECT 57.07 17.295 57.295 17.42 ;
      RECT 57.08 16.585 57.295 16.715 ;
      RECT 56.905 15.74 57.235 16.665 ;
      RECT 56.075 17.335 56.405 17.86 ;
      RECT 56.205 16.835 56.405 17.86 ;
      RECT 56.205 16.835 56.955 17.165 ;
      RECT 56.205 15.695 56.395 17.86 ;
      RECT 55.5 16.255 56.395 16.63 ;
      RECT 56.055 15.695 56.395 16.63 ;
      RECT 56.445 19.655 56.775 20.58 ;
      RECT 56.665 18.9 56.835 19.735 ;
      RECT 56.62 19.605 56.835 19.735 ;
      RECT 56.61 18.9 56.835 19.025 ;
      RECT 56.455 18.465 56.785 18.985 ;
      RECT 56.445 25.095 56.775 26.02 ;
      RECT 56.665 24.34 56.835 25.175 ;
      RECT 56.62 25.045 56.835 25.175 ;
      RECT 56.61 24.34 56.835 24.465 ;
      RECT 56.455 23.905 56.785 24.425 ;
      RECT 55.595 19.69 55.935 20.625 ;
      RECT 55.745 18.46 55.935 20.625 ;
      RECT 55.04 19.69 55.935 20.065 ;
      RECT 55.745 19.155 56.495 19.485 ;
      RECT 55.745 18.46 55.945 19.485 ;
      RECT 55.615 18.46 55.945 18.985 ;
      RECT 55.595 25.13 55.935 26.065 ;
      RECT 55.745 23.9 55.935 26.065 ;
      RECT 55.04 25.13 55.935 25.505 ;
      RECT 55.745 24.595 56.495 24.925 ;
      RECT 55.745 23.9 55.945 24.925 ;
      RECT 55.615 23.9 55.945 24.425 ;
      RECT 55.905 22.565 56.37 22.895 ;
      RECT 56.05 21.605 56.37 22.895 ;
      RECT 54.545 17.625 55.33 17.795 ;
      RECT 55.16 15.825 55.33 17.795 ;
      RECT 55.16 16.835 56.035 17.165 ;
      RECT 54.445 15.825 55.33 15.995 ;
      RECT 55.535 33.655 55.865 34.175 ;
      RECT 55.745 32.905 55.915 33.74 ;
      RECT 55.69 33.615 55.915 33.74 ;
      RECT 55.7 32.905 55.915 33.035 ;
      RECT 55.525 32.06 55.855 32.985 ;
      RECT 55.35 23.065 55.755 23.235 ;
      RECT 55.35 21.135 55.52 23.235 ;
      RECT 54.69 22.535 55.52 22.835 ;
      RECT 54.69 22.505 54.89 22.835 ;
      RECT 55.35 21.135 55.6 21.465 ;
      RECT 53.985 20.325 54.87 20.495 ;
      RECT 54.7 18.525 54.87 20.495 ;
      RECT 54.7 19.155 55.575 19.485 ;
      RECT 54.085 18.525 54.87 18.695 ;
      RECT 53.985 25.765 54.87 25.935 ;
      RECT 54.7 23.965 54.87 25.935 ;
      RECT 54.7 24.595 55.575 24.925 ;
      RECT 54.085 23.965 54.87 24.135 ;
      RECT 54.695 33.655 55.025 34.18 ;
      RECT 54.825 33.155 55.025 34.18 ;
      RECT 54.825 33.155 55.575 33.485 ;
      RECT 54.825 32.015 55.015 34.18 ;
      RECT 54.12 32.575 55.015 32.95 ;
      RECT 54.675 32.015 55.015 32.95 ;
      RECT 55.065 35.975 55.395 36.9 ;
      RECT 55.285 35.22 55.455 36.055 ;
      RECT 55.24 35.925 55.455 36.055 ;
      RECT 55.23 35.22 55.455 35.345 ;
      RECT 55.075 34.785 55.405 35.305 ;
      RECT 53.805 23.065 54.48 23.235 ;
      RECT 54.31 22.115 54.48 23.235 ;
      RECT 55.01 22.025 55.18 22.355 ;
      RECT 54.31 22.115 55.18 22.285 ;
      RECT 54.67 22.025 55.18 22.285 ;
      RECT 54.67 21.24 54.84 22.285 ;
      RECT 53.735 21.24 54.84 21.41 ;
      RECT 54.215 36.01 54.555 36.945 ;
      RECT 54.365 34.78 54.555 36.945 ;
      RECT 53.66 36.01 54.555 36.385 ;
      RECT 54.365 35.475 55.115 35.805 ;
      RECT 54.365 34.78 54.565 35.805 ;
      RECT 54.235 34.78 54.565 35.305 ;
      RECT 54.525 17.125 54.99 17.455 ;
      RECT 54.67 16.165 54.99 17.455 ;
      RECT 53.165 33.945 53.95 34.115 ;
      RECT 53.78 32.145 53.95 34.115 ;
      RECT 53.78 33.155 54.655 33.485 ;
      RECT 53.065 32.145 53.95 32.315 ;
      RECT 54.21 18.865 54.53 20.155 ;
      RECT 54.065 18.865 54.53 19.195 ;
      RECT 54.21 24.305 54.53 25.595 ;
      RECT 54.065 24.305 54.53 24.635 ;
      RECT 53.615 22.645 54.14 22.865 ;
      RECT 53.97 21.58 54.14 22.865 ;
      RECT 53.97 21.58 54.5 21.945 ;
      RECT 53.97 17.625 54.375 17.795 ;
      RECT 53.97 15.695 54.14 17.795 ;
      RECT 53.31 17.095 54.14 17.395 ;
      RECT 53.31 17.065 53.51 17.395 ;
      RECT 53.97 15.695 54.22 16.025 ;
      RECT 52.605 36.645 53.49 36.815 ;
      RECT 53.32 34.845 53.49 36.815 ;
      RECT 53.32 35.475 54.195 35.805 ;
      RECT 52.705 34.845 53.49 35.015 ;
      RECT 53.8 14.515 54.055 15.185 ;
      RECT 53.885 12.975 54.055 15.185 ;
      RECT 53.87 12.975 54.055 13.385 ;
      RECT 53.8 12.975 54.055 13.305 ;
      RECT 53.51 20.295 53.76 20.625 ;
      RECT 53.51 18.525 53.68 20.625 ;
      RECT 52.85 18.925 53.05 19.255 ;
      RECT 52.85 18.925 53.68 19.225 ;
      RECT 53.51 18.525 53.915 18.695 ;
      RECT 53.51 25.735 53.76 26.065 ;
      RECT 53.51 23.965 53.68 26.065 ;
      RECT 52.85 24.365 53.05 24.695 ;
      RECT 52.85 24.365 53.68 24.665 ;
      RECT 53.51 23.965 53.915 24.135 ;
      RECT 52.425 17.625 53.1 17.795 ;
      RECT 52.93 16.675 53.1 17.795 ;
      RECT 53.63 16.585 53.8 16.915 ;
      RECT 52.93 16.675 53.8 16.845 ;
      RECT 53.29 16.585 53.8 16.845 ;
      RECT 53.29 15.8 53.46 16.845 ;
      RECT 52.355 15.8 53.46 15.97 ;
      RECT 50.655 14.175 50.825 15.185 ;
      RECT 50.655 14.175 53.715 14.345 ;
      RECT 53.545 13.455 53.715 14.345 ;
      RECT 52.915 13.455 53.715 13.625 ;
      RECT 50.655 13.455 51.72 13.625 ;
      RECT 51.55 12.975 51.72 13.625 ;
      RECT 52.915 12.975 53.085 13.625 ;
      RECT 50.655 12.975 50.825 13.625 ;
      RECT 51.55 12.975 53.085 13.225 ;
      RECT 53.275 23.065 53.61 23.235 ;
      RECT 53.275 22.795 53.445 23.235 ;
      RECT 53.22 21.56 53.39 22.925 ;
      RECT 53.275 21.135 53.525 21.69 ;
      RECT 53.145 33.445 53.61 33.775 ;
      RECT 53.29 32.485 53.61 33.775 ;
      RECT 51.895 20.35 53 20.52 ;
      RECT 52.83 19.475 53 20.52 ;
      RECT 52.83 19.475 53.34 19.735 ;
      RECT 53.17 19.405 53.34 19.735 ;
      RECT 52.47 19.475 53.34 19.645 ;
      RECT 52.47 18.525 52.64 19.645 ;
      RECT 51.965 18.525 52.64 18.695 ;
      RECT 51.895 25.79 53 25.96 ;
      RECT 52.83 24.915 53 25.96 ;
      RECT 52.83 24.915 53.34 25.175 ;
      RECT 53.17 24.845 53.34 25.175 ;
      RECT 52.47 24.915 53.34 25.085 ;
      RECT 52.47 23.965 52.64 25.085 ;
      RECT 51.965 23.965 52.64 24.135 ;
      RECT 52.95 13.825 53.325 13.995 ;
      RECT 52.95 13.795 53.315 13.995 ;
      RECT 52.83 35.185 53.15 36.475 ;
      RECT 52.685 35.185 53.15 35.515 ;
      RECT 52.88 14.515 53.13 15.185 ;
      RECT 51.495 14.515 51.725 14.845 ;
      RECT 51.495 14.515 53.13 14.755 ;
      RECT 52.235 17.205 52.76 17.425 ;
      RECT 52.59 16.14 52.76 17.425 ;
      RECT 52.59 16.14 53.12 16.505 ;
      RECT 52.59 33.945 52.995 34.115 ;
      RECT 52.59 32.015 52.76 34.115 ;
      RECT 51.93 33.415 52.76 33.715 ;
      RECT 51.93 33.385 52.13 33.715 ;
      RECT 52.59 32.015 52.84 32.345 ;
      RECT 52.45 13.795 52.78 13.995 ;
      RECT 52.45 13.395 52.735 13.995 ;
      RECT 52.13 19.815 52.66 20.18 ;
      RECT 52.13 18.895 52.3 20.18 ;
      RECT 51.775 18.895 52.3 19.115 ;
      RECT 52.13 25.255 52.66 25.62 ;
      RECT 52.13 24.335 52.3 25.62 ;
      RECT 51.775 24.335 52.3 24.555 ;
      RECT 52.13 36.615 52.38 36.945 ;
      RECT 52.13 34.845 52.3 36.945 ;
      RECT 51.47 35.245 51.67 35.575 ;
      RECT 51.47 35.245 52.3 35.545 ;
      RECT 52.13 34.845 52.535 35.015 ;
      RECT 51.045 33.945 51.72 34.115 ;
      RECT 51.55 32.995 51.72 34.115 ;
      RECT 52.25 32.905 52.42 33.235 ;
      RECT 51.55 32.995 52.42 33.165 ;
      RECT 51.91 32.905 52.42 33.165 ;
      RECT 51.91 32.12 52.08 33.165 ;
      RECT 50.975 32.12 52.08 32.29 ;
      RECT 51.575 22.795 51.745 23.255 ;
      RECT 51.575 22.795 52.24 22.965 ;
      RECT 52.01 21.635 52.24 22.965 ;
      RECT 51.575 21.635 52.24 21.805 ;
      RECT 51.575 21.135 51.745 21.805 ;
      RECT 51.895 17.625 52.23 17.795 ;
      RECT 51.895 17.355 52.065 17.795 ;
      RECT 51.84 16.12 52.01 17.485 ;
      RECT 51.895 15.695 52.145 16.25 ;
      RECT 51.705 13.795 52.18 13.995 ;
      RECT 51.9 13.395 52.18 13.995 ;
      RECT 50.995 15.015 52.165 15.185 ;
      RECT 51.835 14.975 52.165 15.185 ;
      RECT 50.995 14.515 51.325 15.185 ;
      RECT 50.515 36.67 51.62 36.84 ;
      RECT 51.45 35.795 51.62 36.84 ;
      RECT 51.45 35.795 51.96 36.055 ;
      RECT 51.79 35.725 51.96 36.055 ;
      RECT 51.09 35.795 51.96 35.965 ;
      RECT 51.09 34.845 51.26 35.965 ;
      RECT 50.585 34.845 51.26 35.015 ;
      RECT 51.435 20.07 51.685 20.625 ;
      RECT 51.38 18.835 51.55 20.2 ;
      RECT 51.435 18.525 51.605 18.965 ;
      RECT 51.435 18.525 51.77 18.695 ;
      RECT 51.435 25.51 51.685 26.065 ;
      RECT 51.38 24.275 51.55 25.64 ;
      RECT 51.435 23.965 51.605 24.405 ;
      RECT 51.435 23.965 51.77 24.135 ;
      RECT 47.895 11.815 48.065 12.465 ;
      RECT 48.735 11.815 48.905 12.46 ;
      RECT 47.895 11.815 49.315 11.985 ;
      RECT 49.14 11.105 49.315 11.985 ;
      RECT 49.14 11.475 51.765 11.645 ;
      RECT 47.815 11.105 49.315 11.275 ;
      RECT 48.655 10.255 48.985 11.275 ;
      RECT 47.815 10.255 48.145 11.275 ;
      RECT 50.855 33.525 51.38 33.745 ;
      RECT 51.21 32.46 51.38 33.745 ;
      RECT 51.21 32.46 51.74 32.825 ;
      RECT 50.75 36.135 51.28 36.5 ;
      RECT 50.75 35.215 50.92 36.5 ;
      RECT 50.395 35.215 50.92 35.435 ;
      RECT 50.195 17.355 50.365 17.815 ;
      RECT 50.195 17.355 50.86 17.525 ;
      RECT 50.63 16.195 50.86 17.525 ;
      RECT 50.195 16.195 50.86 16.365 ;
      RECT 50.195 15.695 50.365 16.365 ;
      RECT 50.515 33.945 50.85 34.115 ;
      RECT 50.515 33.675 50.685 34.115 ;
      RECT 50.46 32.44 50.63 33.805 ;
      RECT 50.515 32.015 50.765 32.57 ;
      RECT 49.735 19.955 49.905 20.625 ;
      RECT 49.735 19.955 50.4 20.125 ;
      RECT 50.17 18.795 50.4 20.125 ;
      RECT 49.735 18.795 50.4 18.965 ;
      RECT 49.735 18.505 49.905 18.965 ;
      RECT 49.735 25.395 49.905 26.065 ;
      RECT 49.735 25.395 50.4 25.565 ;
      RECT 50.17 24.235 50.4 25.565 ;
      RECT 49.735 24.235 50.4 24.405 ;
      RECT 49.735 23.945 49.905 24.405 ;
      RECT 50.055 36.39 50.305 36.945 ;
      RECT 50 35.155 50.17 36.52 ;
      RECT 50.055 34.845 50.225 35.285 ;
      RECT 50.055 34.845 50.39 35.015 ;
      RECT 48.815 33.675 48.985 34.135 ;
      RECT 48.815 33.675 49.48 33.845 ;
      RECT 49.25 32.515 49.48 33.845 ;
      RECT 48.815 32.515 49.48 32.685 ;
      RECT 48.815 32.015 48.985 32.685 ;
      RECT 49.2 23.015 49.455 23.345 ;
      RECT 49.285 21.135 49.455 23.345 ;
      RECT 49.245 23.005 49.455 23.345 ;
      RECT 49.27 22.935 49.455 23.345 ;
      RECT 49.2 21.135 49.455 21.805 ;
      RECT 49.2 28.455 49.455 28.785 ;
      RECT 49.285 26.575 49.455 28.785 ;
      RECT 49.245 28.445 49.455 28.785 ;
      RECT 49.27 28.375 49.455 28.785 ;
      RECT 49.2 26.575 49.455 27.245 ;
      RECT 49.2 30.835 49.455 31.505 ;
      RECT 49.285 29.295 49.455 31.505 ;
      RECT 49.27 29.295 49.455 29.705 ;
      RECT 49.2 29.295 49.455 29.625 ;
      RECT 46.95 23.095 48.485 23.345 ;
      RECT 48.315 22.695 48.485 23.345 ;
      RECT 46.055 22.695 46.225 23.345 ;
      RECT 46.95 22.695 47.12 23.345 ;
      RECT 48.315 22.695 49.115 22.865 ;
      RECT 48.945 21.975 49.115 22.865 ;
      RECT 46.055 22.695 47.12 22.865 ;
      RECT 46.055 21.975 49.115 22.145 ;
      RECT 46.055 21.135 46.225 22.145 ;
      RECT 46.95 28.535 48.485 28.785 ;
      RECT 48.315 28.135 48.485 28.785 ;
      RECT 46.055 28.135 46.225 28.785 ;
      RECT 46.95 28.135 47.12 28.785 ;
      RECT 48.315 28.135 49.115 28.305 ;
      RECT 48.945 27.415 49.115 28.305 ;
      RECT 46.055 28.135 47.12 28.305 ;
      RECT 46.055 27.415 49.115 27.585 ;
      RECT 46.055 26.575 46.225 27.585 ;
      RECT 46.055 30.495 46.225 31.505 ;
      RECT 46.055 30.495 49.115 30.665 ;
      RECT 48.945 29.775 49.115 30.665 ;
      RECT 48.315 29.775 49.115 29.945 ;
      RECT 46.055 29.775 47.12 29.945 ;
      RECT 46.95 29.295 47.12 29.945 ;
      RECT 48.315 29.295 48.485 29.945 ;
      RECT 46.055 29.295 46.225 29.945 ;
      RECT 46.95 29.295 48.485 29.545 ;
      RECT 48.355 36.275 48.525 36.945 ;
      RECT 48.355 36.275 49.02 36.445 ;
      RECT 48.79 35.115 49.02 36.445 ;
      RECT 48.355 35.115 49.02 35.285 ;
      RECT 48.355 34.825 48.525 35.285 ;
      RECT 48.35 22.325 48.715 22.525 ;
      RECT 48.35 22.325 48.725 22.495 ;
      RECT 48.35 27.765 48.715 27.965 ;
      RECT 48.35 27.765 48.725 27.935 ;
      RECT 48.35 30.145 48.725 30.315 ;
      RECT 48.35 30.115 48.715 30.315 ;
      RECT 46.895 21.565 48.53 21.805 ;
      RECT 48.28 21.135 48.53 21.805 ;
      RECT 46.895 21.475 47.125 21.805 ;
      RECT 46.895 27.005 48.53 27.245 ;
      RECT 48.28 26.575 48.53 27.245 ;
      RECT 46.895 26.915 47.125 27.245 ;
      RECT 48.28 30.835 48.53 31.505 ;
      RECT 46.895 30.835 47.125 31.165 ;
      RECT 46.895 30.835 48.53 31.075 ;
      RECT 47.85 22.325 48.135 22.925 ;
      RECT 47.85 22.325 48.18 22.525 ;
      RECT 47.85 27.765 48.135 28.365 ;
      RECT 47.85 27.765 48.18 27.965 ;
      RECT 47.85 30.115 48.18 30.315 ;
      RECT 47.85 29.715 48.135 30.315 ;
      RECT 47.82 17.575 48.075 17.905 ;
      RECT 47.905 15.695 48.075 17.905 ;
      RECT 47.865 17.565 48.075 17.905 ;
      RECT 47.89 17.495 48.075 17.905 ;
      RECT 47.82 15.695 48.075 16.365 ;
      RECT 45.57 17.655 47.105 17.905 ;
      RECT 46.935 17.255 47.105 17.905 ;
      RECT 44.675 17.255 44.845 17.905 ;
      RECT 45.57 17.255 45.74 17.905 ;
      RECT 46.935 17.255 47.735 17.425 ;
      RECT 47.565 16.535 47.735 17.425 ;
      RECT 44.675 17.255 45.74 17.425 ;
      RECT 44.675 16.535 47.735 16.705 ;
      RECT 44.675 15.695 44.845 16.705 ;
      RECT 47.355 14.215 47.63 15.185 ;
      RECT 47.46 13.135 47.63 15.185 ;
      RECT 47.355 13.135 47.63 13.48 ;
      RECT 47.3 22.325 47.58 22.925 ;
      RECT 47.105 22.325 47.58 22.525 ;
      RECT 47.3 27.765 47.58 28.365 ;
      RECT 47.105 27.765 47.58 27.965 ;
      RECT 47.105 30.115 47.58 30.315 ;
      RECT 47.3 29.715 47.58 30.315 ;
      RECT 46.395 21.135 46.725 21.805 ;
      RECT 47.235 21.135 47.565 21.345 ;
      RECT 46.395 21.135 47.565 21.305 ;
      RECT 46.395 26.575 46.725 27.245 ;
      RECT 47.235 26.575 47.565 26.785 ;
      RECT 46.395 26.575 47.565 26.745 ;
      RECT 46.395 31.335 47.565 31.505 ;
      RECT 47.235 31.295 47.565 31.505 ;
      RECT 46.395 30.835 46.725 31.505 ;
      RECT 46.97 16.885 47.335 17.085 ;
      RECT 46.97 16.885 47.345 17.055 ;
      RECT 45.525 14.505 46.695 14.675 ;
      RECT 46.525 14.215 46.695 14.675 ;
      RECT 45.525 14.215 45.85 14.675 ;
      RECT 46.525 14.215 47.185 14.385 ;
      RECT 47.015 13.375 47.185 14.385 ;
      RECT 47.015 13.715 47.29 14.045 ;
      RECT 45.52 13.375 47.185 13.545 ;
      RECT 46.445 13.025 46.615 13.545 ;
      RECT 45.52 13.025 45.775 13.545 ;
      RECT 45.515 16.125 47.15 16.365 ;
      RECT 46.9 15.695 47.15 16.365 ;
      RECT 45.515 16.035 45.745 16.365 ;
      RECT 46.02 13.715 46.215 14.335 ;
      RECT 46.02 13.715 46.845 14.045 ;
      RECT 46.47 16.885 46.755 17.485 ;
      RECT 46.47 16.885 46.8 17.085 ;
      RECT 45.92 16.885 46.2 17.485 ;
      RECT 45.725 16.885 46.2 17.085 ;
      RECT 45.015 15.695 45.345 16.365 ;
      RECT 45.855 15.695 46.185 15.905 ;
      RECT 45.015 15.695 46.185 15.865 ;
      RECT 40.935 17.255 41.105 17.905 ;
      RECT 40.095 17.255 40.265 17.9 ;
      RECT 39.685 17.255 41.105 17.425 ;
      RECT 39.685 16.545 39.86 17.425 ;
      RECT 37.235 16.915 39.86 17.085 ;
      RECT 39.685 16.545 41.185 16.715 ;
      RECT 40.855 15.695 41.185 16.715 ;
      RECT 40.015 15.695 40.345 16.715 ;
      RECT 40.475 28.135 40.645 28.785 ;
      RECT 39.635 28.135 39.805 28.78 ;
      RECT 39.225 28.135 40.645 28.305 ;
      RECT 39.225 27.425 39.4 28.305 ;
      RECT 36.775 27.795 39.4 27.965 ;
      RECT 39.225 27.425 40.725 27.595 ;
      RECT 40.395 26.575 40.725 27.595 ;
      RECT 39.555 26.575 39.885 27.595 ;
      RECT 37.635 14.165 37.965 15.185 ;
      RECT 36.795 14.165 37.125 15.185 ;
      RECT 36.465 14.165 37.965 14.335 ;
      RECT 36.465 13.455 36.64 14.335 ;
      RECT 34.015 13.795 36.64 13.965 ;
      RECT 36.465 13.455 37.885 13.625 ;
      RECT 37.715 12.975 37.885 13.625 ;
      RECT 36.875 12.98 37.045 13.625 ;
      RECT 29.955 11.815 30.125 12.465 ;
      RECT 30.795 11.815 30.965 12.46 ;
      RECT 29.955 11.815 31.375 11.985 ;
      RECT 31.2 11.105 31.375 11.985 ;
      RECT 31.2 11.475 33.825 11.645 ;
      RECT 29.875 11.105 31.375 11.275 ;
      RECT 30.715 10.255 31.045 11.275 ;
      RECT 29.875 10.255 30.205 11.275 ;
      RECT 29.955 17.255 30.125 17.905 ;
      RECT 30.795 17.255 30.965 17.9 ;
      RECT 29.955 17.255 31.375 17.425 ;
      RECT 31.2 16.545 31.375 17.425 ;
      RECT 31.2 16.915 33.825 17.085 ;
      RECT 29.875 16.545 31.375 16.715 ;
      RECT 30.715 15.695 31.045 16.715 ;
      RECT 29.875 15.695 30.205 16.715 ;
      RECT 21.975 25.045 22.305 26.065 ;
      RECT 21.135 25.045 21.465 26.065 ;
      RECT 21.135 25.045 22.635 25.215 ;
      RECT 22.46 24.335 22.635 25.215 ;
      RECT 22.46 24.675 25.085 24.845 ;
      RECT 21.215 24.335 22.635 24.505 ;
      RECT 22.055 23.86 22.225 24.505 ;
      RECT 21.215 23.855 21.385 24.505 ;
      RECT 20.135 14.165 20.465 15.185 ;
      RECT 19.295 14.165 19.625 15.185 ;
      RECT 19.295 14.165 20.795 14.335 ;
      RECT 20.62 13.455 20.795 14.335 ;
      RECT 20.62 13.795 23.245 13.965 ;
      RECT 19.375 13.455 20.795 13.625 ;
      RECT 20.215 12.98 20.385 13.625 ;
      RECT 19.375 12.975 19.545 13.625 ;
      RECT 19.375 17.255 19.545 17.905 ;
      RECT 20.215 17.255 20.385 17.9 ;
      RECT 19.375 17.255 20.795 17.425 ;
      RECT 20.62 16.545 20.795 17.425 ;
      RECT 20.62 16.915 23.245 17.085 ;
      RECT 19.295 16.545 20.795 16.715 ;
      RECT 20.135 15.695 20.465 16.715 ;
      RECT 19.295 15.695 19.625 16.715 ;
      RECT 189.485 10.265 189.775 11.25 ;
      RECT 189.485 11.91 189.775 12.455 ;
      RECT 189.485 12.985 189.775 13.53 ;
      RECT 189.485 14.19 189.775 15.175 ;
      RECT 189.485 15.705 189.775 16.69 ;
      RECT 189.485 17.35 189.775 17.895 ;
      RECT 189.485 18.425 189.775 18.97 ;
      RECT 189.485 19.63 189.775 20.615 ;
      RECT 189.485 21.145 189.775 22.13 ;
      RECT 189.485 22.79 189.775 23.335 ;
      RECT 189.485 23.865 189.775 24.41 ;
      RECT 189.485 25.07 189.775 26.055 ;
      RECT 189.485 26.585 189.775 27.57 ;
      RECT 189.485 28.23 189.775 28.775 ;
      RECT 189.485 29.305 189.775 29.85 ;
      RECT 189.485 30.51 189.775 31.495 ;
      RECT 189.485 32.025 189.775 33.01 ;
      RECT 189.485 33.67 189.775 34.215 ;
      RECT 189.485 34.745 189.775 35.29 ;
      RECT 189.485 35.95 189.775 36.935 ;
      RECT 189.485 37.465 189.775 38.45 ;
      RECT 189.485 39.11 189.775 39.655 ;
      RECT 189.485 40.185 189.775 40.73 ;
      RECT 189.485 41.39 189.775 42.375 ;
      RECT 189.485 42.905 189.775 43.89 ;
      RECT 189.485 44.55 189.775 45.095 ;
      RECT 189.485 45.625 189.775 46.17 ;
      RECT 189.485 46.83 189.775 47.815 ;
      RECT 189.485 48.345 189.775 49.33 ;
      RECT 189.485 49.99 189.775 50.535 ;
      RECT 189.485 51.065 189.775 51.61 ;
      RECT 189.485 52.27 189.775 53.255 ;
      RECT 189.485 53.785 189.775 54.77 ;
      RECT 189.485 55.43 189.775 55.975 ;
      RECT 189.485 56.505 189.775 57.05 ;
      RECT 189.485 57.71 189.775 58.695 ;
      RECT 181.27 21.635 181.46 22.355 ;
      RECT 180.34 24.675 181.44 24.875 ;
      RECT 179.14 21.88 179.38 22.475 ;
      RECT 178.35 21.935 178.63 22.885 ;
      RECT 177.12 16.885 178.22 17.085 ;
      RECT 177.995 21.135 178.18 23.255 ;
      RECT 177.07 21.975 177.42 22.625 ;
      RECT 173.45 16.195 173.64 16.915 ;
      RECT 171.525 24.595 171.825 24.925 ;
      RECT 171.32 16.44 171.56 17.035 ;
      RECT 170.53 16.495 170.81 17.445 ;
      RECT 170.175 24.615 170.64 24.925 ;
      RECT 170.175 15.695 170.36 17.815 ;
      RECT 169.77 19.405 169.96 20.125 ;
      RECT 169.25 16.535 169.6 17.185 ;
      RECT 169.255 23.865 169.515 26.055 ;
      RECT 167.64 19.285 167.88 19.88 ;
      RECT 166.85 18.875 167.13 19.825 ;
      RECT 166.55 21.635 166.74 22.355 ;
      RECT 166.495 18.505 166.68 20.625 ;
      RECT 165.57 19.135 165.92 19.785 ;
      RECT 164.42 21.88 164.66 22.475 ;
      RECT 163.32 11.445 164.42 11.645 ;
      RECT 163.63 21.935 163.91 22.885 ;
      RECT 162.4 16.885 163.5 17.085 ;
      RECT 163.275 21.135 163.46 23.255 ;
      RECT 162.345 19.215 162.885 19.775 ;
      RECT 162.35 21.975 162.7 22.625 ;
      RECT 158.14 24.675 158.49 24.885 ;
      RECT 157.81 16.195 158 16.915 ;
      RECT 157.81 21.635 158 22.355 ;
      RECT 157.525 24.675 157.97 24.875 ;
      RECT 157.35 27.765 157.795 27.965 ;
      RECT 157.35 19.405 157.54 20.125 ;
      RECT 156.83 27.755 157.18 27.965 ;
      RECT 155.68 16.44 155.92 17.035 ;
      RECT 155.68 21.88 155.92 22.475 ;
      RECT 155.22 19.285 155.46 19.88 ;
      RECT 154.89 16.495 155.17 17.445 ;
      RECT 154.89 21.935 155.17 22.885 ;
      RECT 154.535 15.695 154.72 17.815 ;
      RECT 154.535 21.135 154.72 23.255 ;
      RECT 154.43 18.875 154.71 19.825 ;
      RECT 154.075 18.505 154.26 20.625 ;
      RECT 153.61 16.535 153.96 17.185 ;
      RECT 153.61 21.975 153.96 22.625 ;
      RECT 153.15 19.135 153.5 19.785 ;
      RECT 151.82 24.675 152.92 24.875 ;
      RECT 148.6 11.445 149.7 11.645 ;
      RECT 143.54 13.795 144.64 13.995 ;
      RECT 143.09 16.885 143.535 17.085 ;
      RECT 143.09 19.235 143.535 19.435 ;
      RECT 142.57 16.875 142.92 17.085 ;
      RECT 142.57 19.235 142.92 19.445 ;
      RECT 141.12 24.675 141.47 24.885 ;
      RECT 141.12 30.115 141.47 30.325 ;
      RECT 140.505 24.675 140.95 24.875 ;
      RECT 140.505 30.115 140.95 30.315 ;
      RECT 139.41 27.075 139.6 27.795 ;
      RECT 138.48 11.445 139.58 11.645 ;
      RECT 138.95 21.635 139.14 22.355 ;
      RECT 137.28 27.32 137.52 27.915 ;
      RECT 137.11 19.405 137.3 20.125 ;
      RECT 136.82 21.88 137.06 22.475 ;
      RECT 136.49 27.375 136.77 28.325 ;
      RECT 136.135 26.575 136.32 28.695 ;
      RECT 136.03 21.935 136.31 22.885 ;
      RECT 135.675 21.135 135.86 23.255 ;
      RECT 135.27 16.885 135.715 17.085 ;
      RECT 135.21 27.415 135.56 28.065 ;
      RECT 134.98 19.285 135.22 19.88 ;
      RECT 134.75 16.875 135.1 17.085 ;
      RECT 134.75 21.975 135.1 22.625 ;
      RECT 134.19 18.875 134.47 19.825 ;
      RECT 132.96 13.795 134.06 13.995 ;
      RECT 133.835 18.505 134.02 20.625 ;
      RECT 132.91 19.135 133.26 19.785 ;
      RECT 128.83 21.635 129.02 22.355 ;
      RECT 128.83 27.075 129.02 27.795 ;
      RECT 126.7 21.88 126.94 22.475 ;
      RECT 126.7 27.32 126.94 27.915 ;
      RECT 126.07 16.885 126.515 17.085 ;
      RECT 125.91 21.935 126.19 22.885 ;
      RECT 125.91 27.375 126.19 28.325 ;
      RECT 125.55 16.875 125.9 17.085 ;
      RECT 125.555 21.135 125.74 23.255 ;
      RECT 125.555 26.575 125.74 28.695 ;
      RECT 124.63 21.975 124.98 22.625 ;
      RECT 124.63 27.415 124.98 28.065 ;
      RECT 122.38 11.445 123.48 11.645 ;
      RECT 122.38 16.885 123.48 17.085 ;
      RECT 122.39 19.405 122.58 20.125 ;
      RECT 122.39 24.845 122.58 25.565 ;
      RECT 120.09 27.765 120.535 27.965 ;
      RECT 120.09 30.115 120.535 30.315 ;
      RECT 120.26 19.285 120.5 19.88 ;
      RECT 120.26 24.725 120.5 25.32 ;
      RECT 119.57 27.755 119.92 27.965 ;
      RECT 119.57 30.115 119.92 30.325 ;
      RECT 119.47 18.875 119.75 19.825 ;
      RECT 119.47 24.315 119.75 25.265 ;
      RECT 119.115 18.505 119.3 20.625 ;
      RECT 119.115 23.945 119.3 26.065 ;
      RECT 118.71 13.795 119.155 13.995 ;
      RECT 118.19 13.795 118.54 14.005 ;
      RECT 118.19 19.135 118.54 19.785 ;
      RECT 118.19 24.575 118.54 25.225 ;
      RECT 114.56 13.795 115.66 13.995 ;
      RECT 114.57 21.635 114.76 22.355 ;
      RECT 113.64 19.235 114.74 19.435 ;
      RECT 113.19 24.675 113.635 24.875 ;
      RECT 112.67 24.675 113.02 24.885 ;
      RECT 112.44 21.88 112.68 22.475 ;
      RECT 111.81 16.885 112.255 17.085 ;
      RECT 111.65 21.935 111.93 22.885 ;
      RECT 111.29 16.875 111.64 17.085 ;
      RECT 111.295 21.135 111.48 23.255 ;
      RECT 110.37 21.975 110.72 22.625 ;
      RECT 103.52 13.795 104.62 13.995 ;
      RECT 103.52 16.885 104.62 17.085 ;
      RECT 99.85 21.635 100.04 22.355 ;
      RECT 97.54 11.445 98.64 11.645 ;
      RECT 97.88 16.875 98.23 17.085 ;
      RECT 98.01 19.405 98.2 20.125 ;
      RECT 97.72 21.88 97.96 22.475 ;
      RECT 97.265 16.885 97.71 17.085 ;
      RECT 96.93 21.935 97.21 22.885 ;
      RECT 96.575 21.135 96.76 23.255 ;
      RECT 95.88 19.285 96.12 19.88 ;
      RECT 95.65 21.975 96 22.625 ;
      RECT 95.25 24.845 95.44 25.565 ;
      RECT 95.09 18.875 95.37 19.825 ;
      RECT 94.735 18.505 94.92 20.625 ;
      RECT 94.33 30.115 94.775 30.315 ;
      RECT 93.81 19.135 94.16 19.785 ;
      RECT 93.81 30.115 94.16 30.325 ;
      RECT 93.41 13.795 93.855 13.995 ;
      RECT 93.12 24.725 93.36 25.32 ;
      RECT 92.89 13.795 93.24 14.005 ;
      RECT 91.56 11.445 92.66 11.645 ;
      RECT 92.33 24.315 92.61 25.265 ;
      RECT 91.975 23.945 92.16 26.065 ;
      RECT 91.05 24.575 91.4 25.225 ;
      RECT 85.13 21.635 85.32 22.355 ;
      RECT 84.54 16.875 84.89 17.085 ;
      RECT 83.925 16.885 84.37 17.085 ;
      RECT 82.82 11.445 83.92 11.645 ;
      RECT 83.29 19.235 83.735 19.435 ;
      RECT 83 21.88 83.24 22.475 ;
      RECT 82.77 19.235 83.12 19.445 ;
      RECT 82.21 21.935 82.49 22.885 ;
      RECT 81.855 21.135 82.04 23.255 ;
      RECT 81.45 24.845 81.64 25.565 ;
      RECT 80.99 30.115 81.435 30.315 ;
      RECT 80.93 21.975 81.28 22.625 ;
      RECT 80.47 30.115 80.82 30.325 ;
      RECT 79.61 19.405 79.8 20.125 ;
      RECT 79.32 24.725 79.56 25.32 ;
      RECT 78.53 24.315 78.81 25.265 ;
      RECT 78.175 23.945 78.36 26.065 ;
      RECT 77.48 19.285 77.72 19.88 ;
      RECT 77.25 24.575 77.6 25.225 ;
      RECT 76.69 18.875 76.97 19.825 ;
      RECT 76.335 18.505 76.52 20.625 ;
      RECT 75.41 19.135 75.76 19.785 ;
      RECT 74.08 11.445 75.18 11.645 ;
      RECT 74.08 16.885 75.18 17.085 ;
      RECT 74.55 30.115 74.995 30.315 ;
      RECT 74.03 30.115 74.38 30.325 ;
      RECT 71.66 16.875 72.01 17.085 ;
      RECT 71.66 19.235 72.01 19.445 ;
      RECT 71.66 27.755 72.01 27.965 ;
      RECT 71.045 16.885 71.49 17.085 ;
      RECT 71.045 19.235 71.49 19.435 ;
      RECT 71.045 27.765 71.49 27.965 ;
      RECT 70.41 21.635 70.6 22.355 ;
      RECT 68.28 21.88 68.52 22.475 ;
      RECT 67.49 21.935 67.77 22.885 ;
      RECT 67.135 21.135 67.32 23.255 ;
      RECT 65.8 13.795 66.9 13.995 ;
      RECT 65.8 24.675 66.9 24.875 ;
      RECT 66.21 21.975 66.56 22.625 ;
      RECT 63.84 13.795 64.19 14.005 ;
      RECT 63.51 16.195 63.7 16.915 ;
      RECT 63.51 19.405 63.7 20.125 ;
      RECT 63.51 27.075 63.7 27.795 ;
      RECT 63.51 30.285 63.7 31.005 ;
      RECT 62.58 11.445 63.68 11.645 ;
      RECT 63.225 13.795 63.67 13.995 ;
      RECT 61.38 16.44 61.62 17.035 ;
      RECT 61.38 19.285 61.62 19.88 ;
      RECT 61.38 27.32 61.62 27.915 ;
      RECT 61.38 30.165 61.62 30.76 ;
      RECT 60.59 16.495 60.87 17.445 ;
      RECT 60.59 18.875 60.87 19.825 ;
      RECT 60.59 27.375 60.87 28.325 ;
      RECT 60.59 29.755 60.87 30.705 ;
      RECT 60.235 15.695 60.42 17.815 ;
      RECT 60.235 18.505 60.42 20.625 ;
      RECT 60.235 26.575 60.42 28.695 ;
      RECT 60.235 29.385 60.42 31.505 ;
      RECT 59.31 16.535 59.66 17.185 ;
      RECT 59.31 19.135 59.66 19.785 ;
      RECT 59.31 27.415 59.66 28.065 ;
      RECT 59.31 30.015 59.66 30.665 ;
      RECT 55.69 21.635 55.88 22.355 ;
      RECT 54.31 16.195 54.5 16.915 ;
      RECT 53.85 19.405 54.04 20.125 ;
      RECT 53.85 24.845 54.04 25.565 ;
      RECT 53.56 21.88 53.8 22.475 ;
      RECT 52.93 32.515 53.12 33.235 ;
      RECT 52.77 21.935 53.05 22.885 ;
      RECT 52.47 35.725 52.66 36.445 ;
      RECT 52.415 21.135 52.6 23.255 ;
      RECT 52.18 16.44 52.42 17.035 ;
      RECT 51.72 19.285 51.96 19.88 ;
      RECT 51.72 24.725 51.96 25.32 ;
      RECT 51.49 21.975 51.84 22.625 ;
      RECT 51.39 16.495 51.67 17.445 ;
      RECT 51.09 13.795 51.535 13.995 ;
      RECT 51.035 15.695 51.22 17.815 ;
      RECT 50.93 18.875 51.21 19.825 ;
      RECT 50.93 24.315 51.21 25.265 ;
      RECT 50.8 32.76 51.04 33.355 ;
      RECT 50.57 13.795 50.92 14.005 ;
      RECT 50.575 18.505 50.76 20.625 ;
      RECT 50.575 23.945 50.76 26.065 ;
      RECT 50.34 35.605 50.58 36.2 ;
      RECT 50.11 16.535 50.46 17.185 ;
      RECT 50.01 32.815 50.29 33.765 ;
      RECT 49.65 19.135 50 19.785 ;
      RECT 49.65 24.575 50 25.225 ;
      RECT 49.655 32.015 49.84 34.135 ;
      RECT 49.55 35.195 49.83 36.145 ;
      RECT 49.195 34.825 49.38 36.945 ;
      RECT 48.73 32.855 49.08 33.505 ;
      RECT 47.86 11.445 48.96 11.645 ;
      RECT 48.27 35.455 48.62 36.105 ;
      RECT 46.49 22.325 46.935 22.525 ;
      RECT 46.49 27.765 46.935 27.965 ;
      RECT 46.49 30.115 46.935 30.315 ;
      RECT 45.505 14.845 46.695 15.135 ;
      RECT 45.97 22.315 46.32 22.525 ;
      RECT 45.97 27.755 46.32 27.965 ;
      RECT 45.97 30.115 46.32 30.325 ;
      RECT 45.505 13.715 45.85 14.045 ;
      RECT 45.11 16.885 45.555 17.085 ;
      RECT 44.59 16.875 44.94 17.085 ;
      RECT 40.04 16.885 41.14 17.085 ;
      RECT 39.58 27.765 40.68 27.965 ;
      RECT 36.82 13.795 37.92 13.995 ;
      RECT 29.92 11.445 31.02 11.645 ;
      RECT 29.92 16.885 31.02 17.085 ;
      RECT 21.18 24.675 22.28 24.875 ;
      RECT 19.34 13.795 20.44 13.995 ;
      RECT 19.34 16.885 20.44 17.085 ;
      RECT 10.085 10.265 10.375 11.25 ;
      RECT 10.085 11.91 10.375 12.455 ;
      RECT 10.085 12.985 10.375 13.53 ;
      RECT 10.085 14.19 10.375 15.175 ;
      RECT 10.085 15.705 10.375 16.69 ;
      RECT 10.085 17.35 10.375 17.895 ;
      RECT 10.085 18.425 10.375 18.97 ;
      RECT 10.085 19.63 10.375 20.615 ;
      RECT 10.085 21.145 10.375 22.13 ;
      RECT 10.085 22.79 10.375 23.335 ;
      RECT 10.085 23.865 10.375 24.41 ;
      RECT 10.085 25.07 10.375 26.055 ;
      RECT 10.085 26.585 10.375 27.57 ;
      RECT 10.085 28.23 10.375 28.775 ;
      RECT 10.085 29.305 10.375 29.85 ;
      RECT 10.085 30.51 10.375 31.495 ;
      RECT 10.085 32.025 10.375 33.01 ;
      RECT 10.085 33.67 10.375 34.215 ;
      RECT 10.085 34.745 10.375 35.29 ;
      RECT 10.085 35.95 10.375 36.935 ;
      RECT 10.085 37.465 10.375 38.45 ;
      RECT 10.085 39.11 10.375 39.655 ;
      RECT 10.085 40.185 10.375 40.73 ;
      RECT 10.085 41.39 10.375 42.375 ;
      RECT 10.085 42.905 10.375 43.89 ;
      RECT 10.085 44.55 10.375 45.095 ;
      RECT 10.085 45.625 10.375 46.17 ;
      RECT 10.085 46.83 10.375 47.815 ;
      RECT 10.085 48.345 10.375 49.33 ;
      RECT 10.085 49.99 10.375 50.535 ;
      RECT 10.085 51.065 10.375 51.61 ;
      RECT 10.085 52.27 10.375 53.255 ;
      RECT 10.085 53.785 10.375 54.77 ;
      RECT 10.085 55.43 10.375 55.975 ;
      RECT 10.085 56.505 10.375 57.05 ;
      RECT 10.085 57.71 10.375 58.695 ;
  END
END DigitalLDOLogic

END LIBRARY
