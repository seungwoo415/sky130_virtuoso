module inverter(
	input din, 
	input VSS, 
	input VDD,  
	output dout 
); 

endmodule 
