module strong_arm(
	input vdd, 
	input input_n, 
	input vss, 
	input input_p, 
	input clock, 
	output output_n, 
	output output_p 
); 

endmodule
