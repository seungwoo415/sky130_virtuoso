* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : strong_arm                                   *
* Netlisted  : Sat Oct 12 13:52:11 2024                     *
* Pegasus Version: 22.14-s007 Tue Jan 31 16:35:56 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 1 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ptap_tile                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ptap_tile 1
** N=1 EP=1 FDC=0
.ends ptap_tile

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: ntap_tile                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt ntap_tile 1
** N=1 EP=1 FDC=0
.ends ntap_tile

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile                             *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1e-05 $X=570 $Y=0 $dt=0
M1 1 3 2 4 nfet_01v8 L=1.5e-07 W=1e-05 $X=1000 $Y=0 $dt=0
.ends two_finger_mos_tile

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_1                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_1 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 nfet_01v8 L=1.5e-07 W=1e-06 $X=570 $Y=0 $dt=0
M1 1 3 2 4 nfet_01v8 L=1.5e-07 W=1e-06 $X=1000 $Y=0 $dt=0
.ends two_finger_mos_tile_1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_2                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_2 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 pfet_01v8 L=1.5e-07 W=1e-06 $X=570 $Y=0 $dt=1
M1 1 3 2 4 pfet_01v8 L=1.5e-07 W=1e-06 $X=1000 $Y=0 $dt=1
.ends two_finger_mos_tile_2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: two_finger_mos_tile_3                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt two_finger_mos_tile_3 1 2 3 4
** N=4 EP=4 FDC=2
M0 2 3 1 4 pfet_01v8 L=1.5e-07 W=4.2e-07 $X=570 $Y=0 $dt=1
M1 1 3 2 4 pfet_01v8 L=1.5e-07 W=4.2e-07 $X=1000 $Y=0 $dt=1
.ends two_finger_mos_tile_3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: strong_arm_half                                 *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt strong_arm_half 1 2 3 4 5 6 7 8 9 10
** N=10 EP=10 FDC=36
X0 4 ptap_tile $T=0 -29160 0 0 $X=-205 $Y=-29310
X1 3 ntap_tile $T=0 0 0 0 $X=-430 $Y=-540
X2 4 4 4 4 two_finger_mos_tile $T=-430 -26460 0 0 $X=-215 $Y=-27695
X3 4 6 1 4 two_finger_mos_tile $T=1290 -26460 0 0 $X=1505 $Y=-27695
X4 4 6 1 4 two_finger_mos_tile $T=3010 -26460 0 0 $X=3225 $Y=-27695
X5 4 4 4 4 two_finger_mos_tile_1 $T=-430 -14040 0 0 $X=-215 $Y=-15275
X6 4 4 4 4 two_finger_mos_tile_1 $T=-430 -10800 0 0 $X=-215 $Y=-12035
X7 6 7 8 4 two_finger_mos_tile_1 $T=1290 -14040 0 0 $X=1505 $Y=-15275
X8 7 2 5 4 two_finger_mos_tile_1 $T=1290 -10800 0 0 $X=1505 $Y=-12035
X9 6 9 10 4 two_finger_mos_tile_1 $T=3010 -14040 0 0 $X=3225 $Y=-15275
X10 9 5 2 4 two_finger_mos_tile_1 $T=3010 -10800 0 0 $X=3225 $Y=-12035
X11 3 3 3 3 two_finger_mos_tile_2 $T=-430 -7560 0 0 $X=-430 $Y=-9180
X12 3 2 5 3 two_finger_mos_tile_2 $T=1290 -7560 0 0 $X=1290 $Y=-9180
X13 3 5 2 3 two_finger_mos_tile_2 $T=3010 -7560 0 0 $X=3010 $Y=-9180
X14 3 3 3 3 two_finger_mos_tile_3 $T=-430 -4320 0 0 $X=-430 $Y=-5940
X15 3 3 3 3 two_finger_mos_tile_3 $T=-430 -1620 0 0 $X=-430 $Y=-3240
X16 3 7 1 3 two_finger_mos_tile_3 $T=1290 -4320 0 0 $X=1290 $Y=-5940
X17 3 2 1 3 two_finger_mos_tile_3 $T=1290 -1620 0 0 $X=1290 $Y=-3240
X18 3 9 1 3 two_finger_mos_tile_3 $T=3010 -4320 0 0 $X=3010 $Y=-5940
X19 3 5 1 3 two_finger_mos_tile_3 $T=3010 -1620 0 0 $X=3010 $Y=-3240
.ends strong_arm_half

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: strong_arm                                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt strong_arm 3 10 4 1 8 5 2
** N=11 EP=7 FDC=72
X0 1 2 3 4 5 6 7 8 9 10 strong_arm_half $T=0 0 0 0 $X=-430 $Y=-29310
X1 1 2 3 4 5 6 7 8 11 10 strong_arm_half $T=9460 0 1 180 $X=4730 $Y=-29310
.ends strong_arm
