* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : rs_latch_new                                 *
* Netlisted  : Sun Jan 12 00:08:25 2025                     *
* Pegasus Version: 22.14-s007 Tue Jan 31 16:35:56 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 1 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_736669032860                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_736669032860 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_736669032860

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_736669032861                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_736669032861 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_736669032861

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_730309971733                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_730309971733 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_730309971733

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_730309971734                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_730309971734 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=0
.ends nfet_01v8_CDNS_730309971734

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_730309971735                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_730309971735 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1.6e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_730309971735

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: polyConn_CDNS_730309971730                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt polyConn_CDNS_730309971730 1
** N=1 EP=1 FDC=0
.ends polyConn_CDNS_730309971730

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_730309971731                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_730309971731 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_730309971731

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: subTap_CDNS_730309971732                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt subTap_CDNS_730309971732 1
** N=1 EP=1 FDC=0
.ends subTap_CDNS_730309971732

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rs_latch_new                                    *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rs_latch_new 7 1 4 5 2 8
** N=8 EP=6 FDC=8
X0 1 L1M1_C_CDNS_736669032860 $T=1035 -1950 0 0 $X=920 $Y=-2115
X1 2 L1M1_C_CDNS_736669032860 $T=1035 3960 0 0 $X=920 $Y=3795
X2 3 L1M1_C_CDNS_736669032860 $T=1465 100 0 0 $X=1350 $Y=-65
X3 1 L1M1_C_CDNS_736669032860 $T=3435 -2000 0 0 $X=3320 $Y=-2165
X4 2 L1M1_C_CDNS_736669032860 $T=3435 4050 0 0 $X=3320 $Y=3885
X5 4 L1M1_C_CDNS_736669032860 $T=3865 2045 0 0 $X=3750 $Y=1880
X6 1 L1M1_C_CDNS_736669032860 $T=6430 -2010 0 0 $X=6315 $Y=-2175
X7 2 L1M1_C_CDNS_736669032860 $T=6430 4075 0 0 $X=6315 $Y=3910
X8 5 L1M1_C_CDNS_736669032860 $T=6860 1595 0 0 $X=6745 $Y=1430
X9 1 L1M1_C_CDNS_736669032860 $T=8840 -1950 0 0 $X=8725 $Y=-2115
X10 2 L1M1_C_CDNS_736669032860 $T=8840 3960 0 0 $X=8725 $Y=3795
X11 6 L1M1_C_CDNS_736669032860 $T=9270 105 0 0 $X=9155 $Y=-60
X12 2 M1M2_C_CDNS_736669032861 $T=-1945 4595 0 0 $X=-2075 $Y=4275
X13 1 M1M2_C_CDNS_736669032861 $T=13505 -2615 0 0 $X=13375 $Y=-2935
X14 2 4 5 pfet_01v8_CDNS_730309971733 $T=3575 2425 0 0 $X=3130 $Y=2245
X15 2 5 4 pfet_01v8_CDNS_730309971733 $T=6570 2425 0 0 $X=6125 $Y=2245
X16 1 3 7 nfet_01v8_CDNS_730309971734 $T=1175 -1445 0 0 $X=910 $Y=-1595
X17 1 4 3 nfet_01v8_CDNS_730309971734 $T=3575 -1455 0 0 $X=3310 $Y=-1605
X18 1 5 6 nfet_01v8_CDNS_730309971734 $T=6570 -1455 0 0 $X=6305 $Y=-1605
X19 1 6 8 nfet_01v8_CDNS_730309971734 $T=8980 -1445 0 0 $X=8715 $Y=-1595
X20 2 3 7 pfet_01v8_CDNS_730309971735 $T=1175 1825 0 0 $X=730 $Y=1645
X21 2 6 8 pfet_01v8_CDNS_730309971735 $T=8980 1825 0 0 $X=8535 $Y=1645
X22 7 polyConn_CDNS_730309971730 $T=640 830 0 0 $X=505 $Y=665
X23 3 polyConn_CDNS_730309971730 $T=3230 100 0 0 $X=3095 $Y=-65
X24 5 polyConn_CDNS_730309971730 $T=4295 1595 0 0 $X=4160 $Y=1430
X25 4 polyConn_CDNS_730309971730 $T=6190 2045 0 0 $X=6055 $Y=1880
X26 6 polyConn_CDNS_730309971730 $T=7500 105 0 0 $X=7365 $Y=-60
X27 8 polyConn_CDNS_730309971730 $T=10025 980 0 0 $X=9890 $Y=815
X28 2 nwellTap_CDNS_730309971731 $T=2460 2925 0 0 $X=2195 $Y=2360
X29 2 nwellTap_CDNS_730309971731 $T=7840 2925 0 0 $X=7575 $Y=2360
X30 1 subTap_CDNS_730309971732 $T=2480 -955 0 0 $X=2365 $Y=-1340
X31 1 subTap_CDNS_730309971732 $T=7880 -970 0 0 $X=7765 $Y=-1355
.ends rs_latch_new
