module pass_transistors( 
	input Vg_0, 
	input Vg_1, 
	input Vg_2, 
	input Vg_3, 
	input Vg_4, 
	input Vg_5, 
	input Vg_6, 
	input Vg_7, 
	input Vg_8, 
	input Vg_9, 
	input Vg_10, 
	input Vg_11, 
	input Vg_12, 
	input Vg_13, 
	input Vg_14, 
	input Vg_15, 
	input Vg_16, 
	input Vg_17, 
	input Vg_18, 
	input Vg_19, 
	input Vg_20, 
	input Vg_21, 
	input Vg_22, 
	input Vg_23, 
	input Vg_24, 
	input Vg_25, 
	input Vg_26, 
	input Vg_27, 
	input Vg_28, 
	input Vg_29, 
	input Vg_30, 
	input Vg_31
	input VDD, 
	output Vout
); 

endmodule 
