module strong_arm (
	input vss,	
	input input_n, 
	input input_p, 
	input clock, 
	input vdd, 	
	output output_n, 
	output output_p,
); 

endmodule

