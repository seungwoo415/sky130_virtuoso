* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : inverter                                     *
* Netlisted  : Sun Jan 12 00:33:19 2025                     *
* Pegasus Version: 22.14-s007 Tue Jan 31 16:35:56 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nfet_01v8) nfet_01v8_rec nSourceDrain(D) nfet(G) nSourceDrain(S) pwell(B)
*.DEVTMPLT 1 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_736670542250                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_736670542250 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_736670542250

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_736670542251                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_736670542251 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_736670542251

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nfet_01v8_CDNS_730310354533                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nfet_01v8_CDNS_730310354533 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 nfet_01v8 L=1.5e-07 W=1e-06 $X=0 $Y=0 $dt=0
.ends nfet_01v8_CDNS_730310354533

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_730310354534                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_730310354534 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=1.5e-07 W=1.6e-06 $X=0 $Y=0 $dt=1
.ends pfet_01v8_CDNS_730310354534

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_730310354531                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_730310354531 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_730310354531

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: subTap_CDNS_730310354532                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt subTap_CDNS_730310354532 1
** N=1 EP=1 FDC=0
.ends subTap_CDNS_730310354532

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: inverter                                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt inverter 3 4 1 2
** N=4 EP=4 FDC=2
X0 1 L1M1_C_CDNS_736670542250 $T=2665 780 0 0 $X=2550 $Y=615
X1 2 L1M1_C_CDNS_736670542250 $T=2665 6690 0 0 $X=2550 $Y=6525
X2 3 L1M1_C_CDNS_736670542250 $T=3095 2830 0 0 $X=2980 $Y=2665
X3 2 M1M2_C_CDNS_736670542251 $T=-710 7295 0 0 $X=-840 $Y=6975
X4 1 M1M2_C_CDNS_736670542251 $T=5890 105 0 0 $X=5760 $Y=-215
X5 1 3 4 nfet_01v8_CDNS_730310354533 $T=2805 1285 0 0 $X=2540 $Y=1135
X6 2 3 4 pfet_01v8_CDNS_730310354534 $T=2805 4555 0 0 $X=2360 $Y=4375
X7 2 nwellTap_CDNS_730310354531 $T=2920 7265 0 0 $X=2475 $Y=6880
X8 1 subTap_CDNS_730310354532 $T=2735 130 0 0 $X=2440 $Y=-75
.ends inverter
