* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : pass_transistors                             *
* Netlisted  : Thu Oct 24 23:04:19 2024                     *
* Pegasus Version: 22.14-s007 Tue Jan 31 16:35:56 PST 2023  *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MP(pfet_01v8) pfet_01v8_rec pSourceDrain(D) pfet(G) pSourceDrain(S) nwell(B)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: polyConn_CDNS_729836244780                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt polyConn_CDNS_729836244780 1
** N=1 EP=1 FDC=0
.ends polyConn_CDNS_729836244780

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: M1M2_C_CDNS_729836244780                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt M1M2_C_CDNS_729836244780 1
** N=1 EP=1 FDC=0
.ends M1M2_C_CDNS_729836244780

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: L1M1_C_CDNS_729836244781                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt L1M1_C_CDNS_729836244781 1
** N=1 EP=1 FDC=0
.ends L1M1_C_CDNS_729836244781

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_729836244781                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_729836244781 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_729836244781

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nwellTap_CDNS_729836244782                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nwellTap_CDNS_729836244782 1
** N=1 EP=1 FDC=0
.ends nwellTap_CDNS_729836244782

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pfet_01v8_CDNS_729836244783                     *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pfet_01v8_CDNS_729836244783 1 2 3
** N=3 EP=3 FDC=1
M0 2 3 1 1 pfet_01v8 L=2.5e-07 W=1.2e-06 $X=0 $Y=0 $dt=0
.ends pfet_01v8_CDNS_729836244783

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1 2 3 4
** N=4 EP=4 FDC=2
X0 3 4 1 pfet_01v8_CDNS_729836244783 $T=445 180 0 0 $X=0 $Y=0
X1 3 4 2 pfet_01v8_CDNS_729836244783 $T=1505 180 0 0 $X=1060 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pass_transistors                                *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pass_transistors 13 26 27 1 14 15 28 2 3 16
+ 29 17 30 4 18 5 31 19 32 6
+ 20 7 33 8 21 34 22 9 10 23
+ 24 11 12 25
** N=35 EP=34 FDC=32
X0 1 polyConn_CDNS_729836244780 $T=2745 10060 0 0 $X=2610 $Y=9895
X1 2 polyConn_CDNS_729836244780 $T=3180 -2295 0 0 $X=3045 $Y=-2460
X2 3 polyConn_CDNS_729836244780 $T=3800 10050 0 0 $X=3665 $Y=9885
X3 4 polyConn_CDNS_729836244780 $T=4240 -2275 0 0 $X=4105 $Y=-2440
X4 5 polyConn_CDNS_729836244780 $T=4860 10060 0 0 $X=4725 $Y=9895
X5 6 polyConn_CDNS_729836244780 $T=5305 -2265 0 0 $X=5170 $Y=-2430
X6 7 polyConn_CDNS_729836244780 $T=5930 10065 0 0 $X=5795 $Y=9900
X7 8 polyConn_CDNS_729836244780 $T=6355 -2270 0 0 $X=6220 $Y=-2435
X8 9 polyConn_CDNS_729836244780 $T=6985 10070 0 0 $X=6850 $Y=9905
X9 10 polyConn_CDNS_729836244780 $T=7415 -2275 0 0 $X=7280 $Y=-2440
X10 11 polyConn_CDNS_729836244780 $T=8045 10070 0 0 $X=7910 $Y=9905
X11 12 polyConn_CDNS_729836244780 $T=8480 -2275 0 0 $X=8345 $Y=-2440
X12 13 polyConn_CDNS_729836244780 $T=9100 10070 0 0 $X=8965 $Y=9905
X13 14 polyConn_CDNS_729836244780 $T=9540 -2285 0 0 $X=9405 $Y=-2450
X14 15 polyConn_CDNS_729836244780 $T=10950 10065 0 0 $X=10815 $Y=9900
X15 16 polyConn_CDNS_729836244780 $T=11155 -2285 0 0 $X=11020 $Y=-2450
X16 17 polyConn_CDNS_729836244780 $T=12010 10075 0 0 $X=11875 $Y=9910
X17 18 polyConn_CDNS_729836244780 $T=12210 -2270 0 0 $X=12075 $Y=-2435
X18 19 polyConn_CDNS_729836244780 $T=13070 10075 0 0 $X=12935 $Y=9910
X19 20 polyConn_CDNS_729836244780 $T=13265 -2265 0 0 $X=13130 $Y=-2430
X20 21 polyConn_CDNS_729836244780 $T=14125 10090 0 0 $X=13990 $Y=9925
X21 22 polyConn_CDNS_729836244780 $T=14320 -2265 0 0 $X=14185 $Y=-2430
X22 23 polyConn_CDNS_729836244780 $T=15175 10080 0 0 $X=15040 $Y=9915
X23 24 polyConn_CDNS_729836244780 $T=15380 -2275 0 0 $X=15245 $Y=-2440
X24 25 polyConn_CDNS_729836244780 $T=16230 10080 0 0 $X=16095 $Y=9915
X25 26 polyConn_CDNS_729836244780 $T=16445 -2270 0 0 $X=16310 $Y=-2435
X26 27 polyConn_CDNS_729836244780 $T=18100 10090 0 0 $X=17965 $Y=9925
X27 28 polyConn_CDNS_729836244780 $T=18115 -2295 0 0 $X=17980 $Y=-2460
X28 29 polyConn_CDNS_729836244780 $T=19155 10080 0 0 $X=19020 $Y=9915
X29 30 polyConn_CDNS_729836244780 $T=19175 -2285 0 0 $X=19040 $Y=-2450
X30 31 polyConn_CDNS_729836244780 $T=20220 10080 0 0 $X=20085 $Y=9915
X31 32 polyConn_CDNS_729836244780 $T=20235 -2290 0 0 $X=20100 $Y=-2455
X32 33 M1M2_C_CDNS_729836244780 $T=485 12610 0 0 $X=355 $Y=12290
X33 33 M1M2_C_CDNS_729836244780 $T=490 285 0 0 $X=360 $Y=-35
X34 34 M1M2_C_CDNS_729836244780 $T=22800 13950 0 0 $X=22670 $Y=13630
X35 34 M1M2_C_CDNS_729836244780 $T=22865 1745 0 0 $X=22735 $Y=1425
X36 33 L1M1_C_CDNS_729836244781 $T=2480 12060 0 0 $X=2365 $Y=11895
X37 33 L1M1_C_CDNS_729836244781 $T=2915 -255 0 0 $X=2800 $Y=-420
X38 34 L1M1_C_CDNS_729836244781 $T=3010 13260 0 0 $X=2895 $Y=13095
X39 34 L1M1_C_CDNS_729836244781 $T=3445 1045 0 0 $X=3330 $Y=880
X40 33 L1M1_C_CDNS_729836244781 $T=3540 12065 0 0 $X=3425 $Y=11900
X41 3 L1M1_C_CDNS_729836244781 $T=3800 9600 0 0 $X=3685 $Y=9435
X42 33 L1M1_C_CDNS_729836244781 $T=3975 -255 0 0 $X=3860 $Y=-420
X43 34 L1M1_C_CDNS_729836244781 $T=4070 13275 0 0 $X=3955 $Y=13110
X44 4 L1M1_C_CDNS_729836244781 $T=4240 -2730 0 0 $X=4125 $Y=-2895
X45 34 L1M1_C_CDNS_729836244781 $T=4505 1055 0 0 $X=4390 $Y=890
X46 33 L1M1_C_CDNS_729836244781 $T=4600 12065 0 0 $X=4485 $Y=11900
X47 5 L1M1_C_CDNS_729836244781 $T=4860 9140 0 0 $X=4745 $Y=8975
X48 33 L1M1_C_CDNS_729836244781 $T=5035 -255 0 0 $X=4920 $Y=-420
X49 34 L1M1_C_CDNS_729836244781 $T=5130 13260 0 0 $X=5015 $Y=13095
X50 6 L1M1_C_CDNS_729836244781 $T=5305 -3175 0 0 $X=5190 $Y=-3340
X51 34 L1M1_C_CDNS_729836244781 $T=5565 1050 0 0 $X=5450 $Y=885
X52 33 L1M1_C_CDNS_729836244781 $T=5660 12080 0 0 $X=5545 $Y=11915
X53 7 L1M1_C_CDNS_729836244781 $T=5930 8685 0 0 $X=5815 $Y=8520
X54 33 L1M1_C_CDNS_729836244781 $T=6090 -255 0 0 $X=5975 $Y=-420
X55 34 L1M1_C_CDNS_729836244781 $T=6190 13265 0 0 $X=6075 $Y=13100
X56 8 L1M1_C_CDNS_729836244781 $T=6355 -3660 0 0 $X=6240 $Y=-3825
X57 34 L1M1_C_CDNS_729836244781 $T=6620 1050 0 0 $X=6505 $Y=885
X58 33 L1M1_C_CDNS_729836244781 $T=6720 12080 0 0 $X=6605 $Y=11915
X59 9 L1M1_C_CDNS_729836244781 $T=6985 8235 0 0 $X=6870 $Y=8070
X60 33 L1M1_C_CDNS_729836244781 $T=7150 -255 0 0 $X=7035 $Y=-420
X61 34 L1M1_C_CDNS_729836244781 $T=7250 13265 0 0 $X=7135 $Y=13100
X62 10 L1M1_C_CDNS_729836244781 $T=7415 -4105 0 0 $X=7300 $Y=-4270
X63 34 L1M1_C_CDNS_729836244781 $T=7680 1050 0 0 $X=7565 $Y=885
X64 33 L1M1_C_CDNS_729836244781 $T=7775 12085 0 0 $X=7660 $Y=11920
X65 11 L1M1_C_CDNS_729836244781 $T=8045 7760 0 0 $X=7930 $Y=7595
X66 33 L1M1_C_CDNS_729836244781 $T=8210 -255 0 0 $X=8095 $Y=-420
X67 34 L1M1_C_CDNS_729836244781 $T=8305 13265 0 0 $X=8190 $Y=13100
X68 12 L1M1_C_CDNS_729836244781 $T=8480 -4575 0 0 $X=8365 $Y=-4740
X69 34 L1M1_C_CDNS_729836244781 $T=8740 1050 0 0 $X=8625 $Y=885
X70 33 L1M1_C_CDNS_729836244781 $T=8830 12085 0 0 $X=8715 $Y=11920
X71 13 L1M1_C_CDNS_729836244781 $T=9100 7300 0 0 $X=8985 $Y=7135
X72 33 L1M1_C_CDNS_729836244781 $T=9270 -250 0 0 $X=9155 $Y=-415
X73 34 L1M1_C_CDNS_729836244781 $T=9360 13265 0 0 $X=9245 $Y=13100
X74 14 L1M1_C_CDNS_729836244781 $T=9540 -5050 0 0 $X=9425 $Y=-5215
X75 34 L1M1_C_CDNS_729836244781 $T=9800 1050 0 0 $X=9685 $Y=885
X76 33 L1M1_C_CDNS_729836244781 $T=10685 12075 0 0 $X=10570 $Y=11910
X77 33 L1M1_C_CDNS_729836244781 $T=10885 -255 0 0 $X=10770 $Y=-420
X78 15 L1M1_C_CDNS_729836244781 $T=10950 6805 0 0 $X=10835 $Y=6640
X79 16 L1M1_C_CDNS_729836244781 $T=11155 -5545 0 0 $X=11040 $Y=-5710
X80 34 L1M1_C_CDNS_729836244781 $T=11215 13255 0 0 $X=11100 $Y=13090
X81 34 L1M1_C_CDNS_729836244781 $T=11415 1050 0 0 $X=11300 $Y=885
X82 33 L1M1_C_CDNS_729836244781 $T=11745 12075 0 0 $X=11630 $Y=11910
X83 33 L1M1_C_CDNS_729836244781 $T=11940 -255 0 0 $X=11825 $Y=-420
X84 17 L1M1_C_CDNS_729836244781 $T=12010 6285 0 0 $X=11895 $Y=6120
X85 18 L1M1_C_CDNS_729836244781 $T=12210 -6055 0 0 $X=12095 $Y=-6220
X86 34 L1M1_C_CDNS_729836244781 $T=12275 13265 0 0 $X=12160 $Y=13100
X87 34 L1M1_C_CDNS_729836244781 $T=12470 1050 0 0 $X=12355 $Y=885
X88 33 L1M1_C_CDNS_729836244781 $T=12800 12075 0 0 $X=12685 $Y=11910
X89 33 L1M1_C_CDNS_729836244781 $T=12995 -255 0 0 $X=12880 $Y=-420
X90 19 L1M1_C_CDNS_729836244781 $T=13070 5735 0 0 $X=12955 $Y=5570
X91 20 L1M1_C_CDNS_729836244781 $T=13265 -6605 0 0 $X=13150 $Y=-6770
X92 34 L1M1_C_CDNS_729836244781 $T=13330 13265 0 0 $X=13215 $Y=13100
X93 34 L1M1_C_CDNS_729836244781 $T=13525 1050 0 0 $X=13410 $Y=885
X94 33 L1M1_C_CDNS_729836244781 $T=13855 12075 0 0 $X=13740 $Y=11910
X95 33 L1M1_C_CDNS_729836244781 $T=14055 -255 0 0 $X=13940 $Y=-420
X96 21 L1M1_C_CDNS_729836244781 $T=14125 5295 0 0 $X=14010 $Y=5130
X97 22 L1M1_C_CDNS_729836244781 $T=14320 -7055 0 0 $X=14205 $Y=-7220
X98 34 L1M1_C_CDNS_729836244781 $T=14385 13265 0 0 $X=14270 $Y=13100
X99 34 L1M1_C_CDNS_729836244781 $T=14585 1050 0 0 $X=14470 $Y=885
X100 33 L1M1_C_CDNS_729836244781 $T=14905 12065 0 0 $X=14790 $Y=11900
X101 33 L1M1_C_CDNS_729836244781 $T=15115 -260 0 0 $X=15000 $Y=-425
X102 23 L1M1_C_CDNS_729836244781 $T=15175 4755 0 0 $X=15060 $Y=4590
X103 24 L1M1_C_CDNS_729836244781 $T=15380 -7595 0 0 $X=15265 $Y=-7760
X104 34 L1M1_C_CDNS_729836244781 $T=15435 13260 0 0 $X=15320 $Y=13095
X105 34 L1M1_C_CDNS_729836244781 $T=15645 1045 0 0 $X=15530 $Y=880
X106 33 L1M1_C_CDNS_729836244781 $T=15965 12075 0 0 $X=15850 $Y=11910
X107 33 L1M1_C_CDNS_729836244781 $T=16175 -260 0 0 $X=16060 $Y=-425
X108 25 L1M1_C_CDNS_729836244781 $T=16230 4185 0 0 $X=16115 $Y=4020
X109 26 L1M1_C_CDNS_729836244781 $T=16445 -8160 0 0 $X=16330 $Y=-8325
X110 34 L1M1_C_CDNS_729836244781 $T=16495 13260 0 0 $X=16380 $Y=13095
X111 34 L1M1_C_CDNS_729836244781 $T=16705 1045 0 0 $X=16590 $Y=880
X112 33 L1M1_C_CDNS_729836244781 $T=17830 12075 0 0 $X=17715 $Y=11910
X113 33 L1M1_C_CDNS_729836244781 $T=17850 -260 0 0 $X=17735 $Y=-425
X114 27 L1M1_C_CDNS_729836244781 $T=18100 3650 0 0 $X=17985 $Y=3485
X115 28 L1M1_C_CDNS_729836244781 $T=18115 -8740 0 0 $X=18000 $Y=-8905
X116 34 L1M1_C_CDNS_729836244781 $T=18360 13255 0 0 $X=18245 $Y=13090
X117 34 L1M1_C_CDNS_729836244781 $T=18380 1020 0 0 $X=18265 $Y=855
X118 33 L1M1_C_CDNS_729836244781 $T=18890 12095 0 0 $X=18775 $Y=11930
X119 33 L1M1_C_CDNS_729836244781 $T=18910 -260 0 0 $X=18795 $Y=-425
X120 29 L1M1_C_CDNS_729836244781 $T=19155 3160 0 0 $X=19040 $Y=2995
X121 30 L1M1_C_CDNS_729836244781 $T=19175 -9235 0 0 $X=19060 $Y=-9400
X122 34 L1M1_C_CDNS_729836244781 $T=19420 13260 0 0 $X=19305 $Y=13095
X123 34 L1M1_C_CDNS_729836244781 $T=19440 1020 0 0 $X=19325 $Y=855
X124 33 L1M1_C_CDNS_729836244781 $T=19950 12080 0 0 $X=19835 $Y=11915
X125 33 L1M1_C_CDNS_729836244781 $T=19965 -260 0 0 $X=19850 $Y=-425
X126 31 L1M1_C_CDNS_729836244781 $T=20220 2685 0 0 $X=20105 $Y=2520
X127 32 L1M1_C_CDNS_729836244781 $T=20235 -9705 0 0 $X=20120 $Y=-9870
X128 34 L1M1_C_CDNS_729836244781 $T=20480 13240 0 0 $X=20365 $Y=13075
X129 34 L1M1_C_CDNS_729836244781 $T=20495 1020 0 0 $X=20380 $Y=855
X130 33 nwellTap_CDNS_729836244781 $T=1780 12560 0 0 $X=1335 $Y=12175
X131 33 nwellTap_CDNS_729836244781 $T=2175 195 0 0 $X=1730 $Y=-190
X132 33 nwellTap_CDNS_729836244781 $T=21155 12545 0 0 $X=20710 $Y=12160
X133 33 nwellTap_CDNS_729836244781 $T=21200 -5 0 0 $X=20755 $Y=-390
X134 33 nwellTap_CDNS_729836244782 $T=10020 11065 0 0 $X=9755 $Y=10500
X135 33 nwellTap_CDNS_729836244782 $T=10390 -1250 0 0 $X=10125 $Y=-1815
X136 33 nwellTap_CDNS_729836244782 $T=17170 11125 0 0 $X=16905 $Y=10560
X137 33 nwellTap_CDNS_729836244782 $T=17300 -1255 0 0 $X=17035 $Y=-1820
X138 33 34 6 pfet_01v8_CDNS_729836244783 $T=5175 -1865 0 0 $X=4730 $Y=-2045
X139 33 34 8 pfet_01v8_CDNS_729836244783 $T=6230 -1865 0 0 $X=5785 $Y=-2045
X140 33 34 9 pfet_01v8_CDNS_729836244783 $T=6860 10485 0 0 $X=6415 $Y=10305
X141 33 34 11 pfet_01v8_CDNS_729836244783 $T=7915 10485 0 0 $X=7470 $Y=10305
X142 33 34 13 pfet_01v8_CDNS_729836244783 $T=8970 10485 0 0 $X=8525 $Y=10305
X143 33 34 14 pfet_01v8_CDNS_729836244783 $T=9410 -1865 0 0 $X=8965 $Y=-2045
X144 33 34 16 pfet_01v8_CDNS_729836244783 $T=11025 -1865 0 0 $X=10580 $Y=-2045
X145 33 34 18 pfet_01v8_CDNS_729836244783 $T=12080 -1865 0 0 $X=11635 $Y=-2045
X146 33 34 19 pfet_01v8_CDNS_729836244783 $T=12940 10485 0 0 $X=12495 $Y=10305
X147 33 34 21 pfet_01v8_CDNS_729836244783 $T=13995 10485 0 0 $X=13550 $Y=10305
X148 33 34 31 pfet_01v8_CDNS_729836244783 $T=20090 10480 0 0 $X=19645 $Y=10300
X149 33 34 32 pfet_01v8_CDNS_729836244783 $T=20105 -1870 0 0 $X=19660 $Y=-2050
X150 1 3 33 34 MASCO__A1 $T=2175 10305 0 0 $X=2175 $Y=10305
X151 2 4 33 34 MASCO__A1 $T=2610 -2045 0 0 $X=2610 $Y=-2045
X152 5 7 33 34 MASCO__A1 $T=4295 10305 0 0 $X=4295 $Y=10305
X153 10 12 33 34 MASCO__A1 $T=6845 -2045 0 0 $X=6845 $Y=-2045
X154 15 17 33 34 MASCO__A1 $T=10380 10305 0 0 $X=10380 $Y=10305
X155 20 22 33 34 MASCO__A1 $T=12690 -2045 0 0 $X=12690 $Y=-2045
X156 23 25 33 34 MASCO__A1 $T=14600 10300 0 0 $X=14600 $Y=10300
X157 24 26 33 34 MASCO__A1 $T=14810 -2050 0 0 $X=14810 $Y=-2050
X158 27 29 33 34 MASCO__A1 $T=17525 10300 0 0 $X=17525 $Y=10300
X159 28 30 33 34 MASCO__A1 $T=17545 -2050 0 0 $X=17545 $Y=-2050
.ends pass_transistors
